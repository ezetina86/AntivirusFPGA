XlxV38EB    5ec7    16d4�� �/��p	�r|��_�K#=5L=#������ӎn�:++  �DY�*�ޟ�Y�N���VڦO��ћ���Wò;��T�ɫ0B�� 	�a�B��+�G%�F��:yob։�:4:��*U�sP���:�%V���8�#$���r�{���I�&�L5|�]��N�3?ݾ��R�f��5@\�t��Y��?^�ʕ)<}&c�m�Nڊl>�Qߊv��H����}�I@$UƟ��i��<8�$RK�s�jlS�	�wڊegX�^8^Gsz�:�~C�$�McdD�����yՇ��~���2w" %�#�MO�f��!	�����5^��"�$e��fx�/Jwc�Gxl,t�z65��yȀ����S��W���M���-V�uPLo g�4)��O�[��IT��n�9o�[�G�tkM�A+��ĕ:�bL�"�R�}T��%-T��әݴ�Uu�:8�'h�J�ܥ�?������T��ͺ	V���p���B��ėd��}pѠчw�\�K>�`�����:�ALϙf�t�#�C)�!e���N1R�Eы]�ʦ֛4���v��4Y�%c;��z��;ڙ�Z��\��)�7��9wky�u*��'8od�l��K9����/��9�^�M/$���dR�?�dHt¯���5�{�X�����"ՆW��Z{h��s!���g{����}�#�9r�)���I�~}-�nP�9avd��!�4?��.Leq��3��,���s�c���e��}�(��Z��`��o�o�68�
�X!A#ң����Z\��7.3-u�O�V:�x�P���^sW	���欿�w?�B�.SI��G$ ɴE�ѥ�x �>Ә��*�.[�ǁn��\��A@-_G�/�g��sz`�����C]�km��
��Lq�
����&�� ���Q��o�V�/�A�y�Yƿ��#���myo@�ٻ�@D8�u�~W�l�m�0��	�E�V��l�_T�g�ф"�T2�q�lYDS��#�T%�g���`/���FsqsTYW5G��v��;Z�b�u�u:dGR�f$%ڈ�vȕ�@.�gޘ/V�*�>���+.��Y�i�Ѓ�ʉ�Tn�Ϫ��Ha�L����.��v��@�fE{��kK��|0�"�xs��+�!D-�Ƕ��˵U����z}Y�̫7����p�Z�ٔ7�����P��I���=��<�pf��R���<,�P���W���1��������WK�d.�"J�;�����f�3�́-y��`_��P쳫'�MT���=�>1��78��I�/cE����+�;@�2��g����GQ��<a:�橡� C?|�1�^��|5�t&�?�wu͵��=����/�{{Z�GJ��\�����-�l��y�a�#H&K.Np&������m�t���g�M͒��%�m��d�:��Ci�b+l�h�)ɧ��I��hA7u����� b ��Sį�K�)Fz bA�
çP�m[c�.^�"�Ќ�|���bT^�#$�;
��og$��V;(��?�k��0�ٌTeXV<���O�W j�J�3/���D��ΰ3��z#!9n9����������7s����mR��.��b%K�\s�Xg�>�ﭥ<�w���#����a/+��z��T����%�|̨�e���*�����ۀy��xaZ\/g(|�:s�4�,��6_I2�8����p"Ш̗�$%f]�3x}&���H����yck[����P�s%����z*��������)�:���R��H'�
/4��n�7��^<��C	Sϋ��d��� ��)���:��Z���4�]}�ç���g����	$RVͶ*�Vd��%�19�$�+u]̺u!��d�k����a���HG=��g�+~|-��N|J,�s�Kt���=o��e(00�8q��;�s���٣v4Ln��RI��O��i�N�>���|Zjoi����<���)v7�)P͖ȏ�l�H��B"oiv/g��x�㙯���:w	�+c:��^��[i5y�~����zN��_R�_���+�fn��������׼���u	��P-P%x.n+�a��mK	��N�����:��J?���������s��(^�֕������ʦ����ȋ�~��ݩ�F�y��� �d���^��b�"4|���Bn��)����h+��~���yF!��>ѵ�
֦�4׆�㣰p��hr�!��.!�z��\,�a�Gy����V�2��{�*/^�|�6�i`��C�4b��`y�y�P���|��SVޡ�	����g=�}��H��3g%⻐��%����'���)��(��:���SNb��4�f�����W���(Y���I��'�C��Q?�gFЙ��+)���j����	��]8͖�ߖ�PHu���W`��S��:)��{�6���ˤv	�*3
�A��)��?�c'>H�d8�o�:a~�+�@4W�M��/�{v�_԰U�#"�����w��&g�.��X�	U����P@��l�.B-@�A���˥3�d�� �ȴ�V��T��~�˂��GK�ݫ�G༪:�)6�@�G�UN�qE\�(�,�-^��e�\�#0d�G�u7
O�
�`�������g�5�J:ή���w�;�臨��(��j�ǳ��+=S��6�5� -j�s���EJkz�Һ���t꯯�1�J�	��F*a�ilq�46{-�a�
��P�;Ĵ}k����f�cZ�b����MH�'[�k�NOc�.
<e��#��հ�vo�&A]�8#c���J�/9>/�����uT����_��gh�ӯ�{�F6���j��,;*������ԇq�Dr��Ý�^��1��QJ����dS˻��R�.\�n$c��n��1�9 ��j_��>��gw]����PEJn�SJ�;
��OrZE� Q����lThԋ�>(�1X����t<�j3>��R��ɣH�$R`��n^9�.�#�D��O��t)?r�n�z�q{6tP��O��c�K� W�rȰ���n�n0#
1Z[�O�#:3Г���!�C/6�n(�C��x�BTV�I2�[#S���0�n+���C+���fD��U�p!�R�
�ݳ��/V��0Bs�A�Z�Z��_[�bc��� gh�Q�A��X|��(h�W�	9K�
!��R����w7.d1���h�����ro�|��O��m��5)Ğ��s��H��7�@�a��VeB���S�U�co<�D��|q������G"(��� ��cX�����S%|��~����G������ܕ������ŝ�������C����; ��p��cVI͵��~�ɶ�GL7ɯ	35�L�9pOĐ�te���1!{�WT���u	b�:*;��uyw�3�[R��p�z�+B�J7<�q��\���V�:Ҧ`�3!-Y��l�%;�ps��:������!gHFk�La�����촴N�k�<�4O��z���/0s���cDBDb�n%�Qz��N�|5��)� E-*%���"�}w)l�t�.r6��������"�8�]�x|����xGO��7�ː,،̒ȸܲv�_�djo}����"6��<�;H����[!Ů�L��^=F2�(w�޽�(_i!�� ��AFϺ
��������*�5a77��g�4�B5OA�����O�FC�;����\��!&��.U�:,=��d��!l�	�j�RJ j]\ϥ��d����)9���j���Q77y^ݚB�Ի�1�	�H[\�5���o>Yj�|A�8"�h'1[�-� �rε�Q;�
/��SN�}줿��ŢA-sZ����>', ��B���/�VeGG;b��<U#����5V�}�d��H��Z����h3yx|��1�g��b�KmM���yY���\�
#.}�x��e��~����L�*;(�)s0��[~�"%�v�� �Cr�7�?)I�F�����M��z����"e3�Ɠe�t%�Õ�-^).�h��W+D#�:J!J�}���j9O�dx}.y�eU����1�{Qaغ�#�uSA��9KP��W��r!�'�V�d �t�ڲs8�գ�A�|�PA����{-a���dPQ�n�6�
�p=��~h�������U�Ё��&�E��@�}3�e;�v��e��ڗ�z.V�:���t7��ΰ�(�����υw��g��F���E�����dx��� �~B��`Z"<�ur�6T
���S�[����eA�6K��
�V�1G�-Y�83�N�ʅ��ۺ�0CU	������6���Ru�Z�3�J�r�B��� �I�`ǜ�u��Vl����G��K+�9h��t� ������=��<v�Wۜ�<:X��j&��4Ke��\&G<g1b��.�F֞� �!R�G�����&U����0�5���  �>�{��m���ZByA�s���JDU��ht�;psc��)kF%�h�o��z���yc!�\��Oy���_ 0|�KY! �c �rN����e蕥��,8,��L\��fb�\H��B ٱ�
v�, ���ë�6���u�)z$ĄK�}$f���̣�i�� [�!�l5O�~��p�$����Q�Q�y���X�yI��c5�]�Eh��Ԯ��7Y	$���}r�㹪��f���k�fx,�mWr�D�(�{"m�x~���E�~ǧlt�6���)����x$;��/��#dxgx������ahW"L�����CU�(�>�D( 0]W�6���a�t���.u���j3����q�Y[�:����w|��������N�t���`[�`fpy��[���o�-7�p���Gik�!���G+x��:�E#����S��o&ҋ����>Q�D�ƣ�vE��3�P~2|1����tKy����5s�q���m�e�`\fC1�"8d����TC-���ܼe�����9��Ñ7�_���[uqiˋ|��*u��^��?�����-Z�pv�R������R98Y^_n_���B�9R�0F�{�T��I2�QL�	Ħ@�	 �r�[u�k$y�{��9�k��_0o��?�Ye�HO(`����,G�5���/�s��� ζp�T����tLǻ������G�2à����t��]s��l���K����UB�����Љ�%&���Y.�!�s�s�<�TB<��ﶛ��MҤ�\�vN��{�tG�;2?hP+Q��4_�s�h@8w0wQ���!�Δ>���� i�f�h��!���[_R2��f���S���r�p�o�M/�	�5c���`����̦B\���f����q�b��'��n�=5̚5`�2��j��:�}��Yu�����n˖7P����A]q�\�����U{��$�l�I���m�F~��A{#��j`v�N�G�f��[�*]&Zk�h���ԙ��>�:2_���A+�� 5���k%!,K�Ʃ�7%Tk��|�⣤	�Ís�\�jkD��1^}�1h#|6��r�r�̴��?���{�}w5tX-W�8 �BZ�^�|5�P���If���j:�X��N�e���@�g˚@G�D_��,��,���#w$���$\�	�a�aH��;��\!��11�h��Z'B\�-{�g���Ǿ;W���q��T�7�y֓�VY�cj9f�qZ�Vfj�O����z1���^�L�&����j�^��%�\w�^9cɶt�}"bC���c���y%j�vu�r���YS�=�-�M�x�:�@@6<uj
@y�9B~�u���j��j͸<����Ȕ0C��\V�ʼY�[i�aQ����,��