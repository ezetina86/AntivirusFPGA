XlxV38EB    1b3d     6e0�y8�	�(�X	��"2i�?:�ERM�`���uN�wm! {L�,U0	����g� ��0���MMo��Z�K�DE܄�1QA�A!�7�}�mg�1��62`�$��-^��-���0]�#��}-���^��I�'��?�~�e���Am@�BĖ؟��M}�t?��A�PU,4�(�r4Tk+�����6�1v�����0�F��p~T��$���9��5�
�Lf��'����xQc�a����#��ǘ6>���Qb|�v��p�(� �Dq޳�@y�j=������5ۙ��*;b`5|���҆�xp��\�G���aMa�y8� o�2݂�4p�j2~�	����)1u]k�,l[�J
Әv9�9�y���q��U$zq��T-�]��3�j�5E� _�n���L�rl�|YW�>D3�{(�q���ƈu�b%`L[���������-1ƖiX0�N�dH�f�ݷ�D�n���Y]��茛�h���!��*�|ֽ/�ʟw+�Ƒ)i'G�0��:Կ�ŀ�Ӄ�p��
���;Ĭـ���\��!Y�_l||�٥�"׵
�w��Pf^ff���W��#VG&�G���ܞf�G��,�UÔS�4o�w��YͶҡ���_g1��th���{�Sg�?	4W���퓽/E�	V��+�4�����tݗ�I��=)<�uO\	i��u�Di\W"`zl^��+�#�%����/� ���^N���偌HW�A�5��q�,�Fcl�7u���GKp�i�oB�R�(���$=e�¸���#����pp\e�֪6�y�
�i�>�Jv*],8���	�^����D��G#q��s39Ξ���tb���>`AK��`nH���1�ܘ��{�����_l�2"�n?�@/�/s_l����ό ����+��*�~�c�t�9��-Z�,fd��ۀ��?fa�����חn���7�&Q��r�I:Yg�y9 �ŧ[m"�7u+M�vP���ꬔv�Mx(s�>Z�<�N��[l栀g9p��f�nL���% ��JJ��o�K�*�W��g�ݫׇ���k9�}W��K�:�彐fr���"����#(���O�����P�Z!��kLoo���b*��X��50�xW���XyR�'�gt{Z��Rx�hj{�y��0�c~Y��72Ԯѳ��[b*�0�)쬭&X3(��|�$S�O��	�B>z� ��%��)F�UYjV[
t͸�1�^�S���se^���QY�r��ݻ�؅j��G/2��`7�dQ?mb��J��˽U��X{��]�|�b�Z$I�S�E�z��W��vr��fP�a�R�PU?����5�"3]�E�/�3�߇=���{Sb���?g1峺��!ݓF�l��Ml�tWMS ��~!]�b��4�4��o#\ن>O��#�x�������9�,F���Ȝ������f@�=�OWU�c�P�'g��ن��DE� klB�w����S�l��
�C� "Z��s=���  �E��j��qU�A�%�qU�������fL��.M��[�_��������-1D1�"����c��ϩ�F���ٙ�hL�������c��/�@.��!���XL,�x��r�@zԄ>��QM�s�([yi�ӛ�Y�V�����.{����0�Q��Ş ,Sƾ��W�M��ZM��D���>����*9�f�j�26I&������v��Y