XlxV38EB    2525     876|�4�֛L�����S�w�X�0O��������F�}X����-��8�|�ClY��@�\y��Y�i�O�LR���Y6R�R�#O��,��s�Ð�.�E�/����)��V��f1������14��sڶ.Vw����� ���~��@}3��d� �)X�C�������%.?>S�\���W� ��A �������w3�}w�Կ~#}��������[UWWz����:���R`�y�v�w�K�?ʓ��c��c���X���Q�Y��D��-;�
/�������v�G�*�����P��D%��ba�&�b��U�_��h$��@�&�6q�=1�=m�*��c��NS�r�@�E�2�&���E�)�E�š:4�E�4 �z��H��%d��_~����ԩ���]�~���v]3�v�Qd��_��\���8�F�@�c��-u��d��܇��x\��,��C ����x���nC�*E���KmC�;͸��ݩW?!Ogx��+*[fZ�2|{��F�87��Z�5YI�D0���A�k��]��W��]bZa�|�_�YU𝨢��:�vH�)QN�kY���I�i`�­ݰ�N�R�� ���#CS,���⭟�����س�.Ay�	���_�� hk����0X�s*�)��l�̍)�*��4���׳��>G��4'��)LS�Z���aL�[:�[K��Y��YR����yCֻ���>-��)�T�2}+�!N�%�������C���w�������:����)�c�v�I��/���1������"�+ۀ��˕D�1a�*4���v.LC�����ϕ�&Eu�m-����n�#��:;0L�^�%i�}�C/&�����v
�)��e��.�a�J
�E#��"\d{�����6�S���D�ORȶ>7 z&�0z9�m�#�5���{17+,��� �V�Cs�����l��n�v��zcYvl�)\��Q�u��X�	�y��3K��_!��ܬ%����6�JqTٿ��G�=>`��x���������V�q�?�DP��0<#��wY��Acoc���(Ҏ���ۆawJ��1V��6�}�S�7t�t|�*[p���14��v���G�d{�DB�ؔbY�84"Nt��ј��?5a�J���6��j9���2�B����]*�+��O����]�C�,J�y�3���QoN�;*A~ ��N�5���Ѫ,L�N��O��ϗ�r��p��Ġ}�]�K �zbOo{i$�\1yV��:��B��o���(�iէ�ǫ����&��i�ClN��BA�S!�?e��N��]�YU�\"�11u���I�2�6���|?�'�@RKڥ{�T ����LFp@o���j2��AD:WF���� � ��j��jH�-��o�U��`
2�=1`��c��6W8��g����6[��uFi^�m5Tǿ��1�~��K.��F
nN;��M#��x�a�J+Ӹ�c;�\����(�I��~��#�C�ԴX�z�Ό��!{-�%k�y/V��RoGB'��Ι��C c�9��YR�Cᅢ�e�(b�6�cn\#!B���G`�j���Nï�R��]�Ip���^�P�	�s�{b�����k��N'��|E���� 3R�#t�%����T`�\ѦH�4��j�����c��:�@l$$qw	��������1������t !�B�gM]�B*�k[S�G'���3���H�b�X�������D\ϣ����E��K�;��=E\ؽF�₶}�� �����w�B�nm�o[~���K9ǚyZ�fjV_fs�y��Z�<��?���[z~�A$�&��p׸��gӊ:j?�WI��h��;vo�9�l���f���=uVң9Ǜ8�Z��Z]����eٽ�������k?�J��+«XCdF��Zt9���z���u�dX�^�
��N���15���aC��!~�W�Y�����_�R� ��{+�%B�� Oœ�L�U=7�D�q8�d��t`��&=����خ��#?�}'Zi�w�k*�58� �J<�-�9��ܢ��ld�7Yq��t�n}9�!N}�(<��H~�$�Ѐ�5�"(��c͖���5�K��̈