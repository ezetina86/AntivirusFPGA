XlxV38EB    2804     c62"vCˈ#�� �8;S�?�����9d#\~����B<Jk0�?�7�M̳�t/ԺBQFΎr7W�Z�<h{�a)o�f�G�U�7L_���n�����_j�`=�~Q,k�:�����e��� b���n���xax �SF�2�J��}��VU�m\���c4�ܛe�q`k�c�j�Q�|��7�i�&�(��g����^9w�ض}9�W�U�Ɋ�0o��y�/���kI��kX�}]��<�#jV�BT{s��VO�S� �|�0=�GPrYx0��G]�n���>r����f�B����& ����_��z�h�-1,�����돲�ӏ��ZɉҬ@e�5j�j��ی\fE�T�W���fhj�_]��,�U��#�IY �I֋B������"�*��:d"�4��48
���������ґ�����A4Q����-Wg��I���5��q��儀u{0&	�\��ٌc�վ�W��0
����[@o��s�E�0�-��KfA�X��j����U^s��׃�j��/�{N�ҽ����R�+847Q��;�����'f�Y�Ց�_���zN�w��=b<A.��B���Q�$/�#2�d�a��awt<��j�}|�o�E��u��eq�m+	U��2���|!����X��}P������;UI��e8���'��5�[fL���Gqz�q
����ѽ8q޷����;������ugR��)�623���a��ַ&C����;�a�?�d#VX
������J
}8&��W��K�U#�3hp�f���x �?¡Y��0�(�����䓽�HP�$��zz���eO^_YU]^��*JNܡ&�)(��Ζ�����~�j!]��8{�P��zS2����$!X	Z'��`���5�Ϟ?@ն��+�J*�̯���H}����=l����C`\Q�N)��SX�*�8�.�xV�g��5�']�p�Ic�#�o�V�(l#<���,	�cA��eP���70|rr�^ŧ�}�*w	y���o�j]���m������/\�7)����7�Ǝ��pgm��
���$�2�aĻ�9 �����ޱjw�2�z����sN�__�n-��H/�l�W�t�*K�{_;�ρ�[9#��=�n�ʯ���n�*���r�y2 <!"$�۠�*��7^�L)�!o���NEsq0�׈x����� ��=� m�� ?���8A�d��z^]{wd���M�+c�L��W��Y�`)���L	�n��z~nd�G�q_e
&��g�l�a/�A_�V�hL�qQn)��^�%�r�D+�%v�#S�miI�>S� ���D�	�����r`��9dS0x�.Bٱ&-i�4�(٠ٺh���[8�Q�$�9�߄����!���Bs��~&��e���)KM�����5q�:�߼��_��b�%�P"��W�a�s�"֬{nRѠu�s��2�;N*Ԛp'Kf`������Z�xa�M���߇����S�W���AVu�	t@�x�?�H�(5�H�`;t����d:3G\���Yy�mWj>�~�Ex��?�b5`+�P��v��|A�]�f�I�N����"��`���]v�8z�;h�4�A{쭮;B�m���蓿M
hsL 0�:^���P�F�5b�h�~��N�l7o����gͻ�y0R�,�F����u�/�>`4B��VB����TnK����h�T�|�ݮ�1]�������G)1��Sy�� ։�(�M'�>��7��@�GO�we���+���������xJc�2���s����6~F\I7=j�"��OU}�NRc~��n`�$��6�C��Rt(k<����('�J���|�f9�ٲ:C�� Gq��jy���+u��������K���z�x�͡;�$ݏ��Z����	�ʃ����\�Hy�#�]��/��u���>���xT�]�kcm�K���X�M��-K��F&��!�~'���u�BJ�b��ߤ�dDP�	���'3��g�fAN�o��v�t9�����@�'���8V;D:��pF �o�-|,��i3�� �~� ���m[#ʥ;O�{l���]�������K��﬇@4���AMu?A�����>ͷ��Rd7smeؘ��D��&�R|O��+%�tnU� �V�z��\q�Y8���-�vu�w�V��>#����Jɬkxr:���?�E֍Ȁ��G�^��M�3��
v؆�z?h
��kT~9e�`BYX)�`ƶ�:{� �9釽by�R��ݨrC�5��a���>�����Y�<�G��)�
�Ræ���F��-�B.�*hJb֌�EMX�.�3]s�9�����0F>�岽^8���O���vG6jϯɖR6��`f�M�� ћ`�y@�C)�Ţ�#�e�yt��d��⛊1��ޚ�D���U�T\�TJ]5�\�U`�|�4�/��Z�+#:�jj�؞�J�������z�fK`�5Q�[A�y�ќ�2?N1�[�&���
��C�?�s0���du�M�$����ʾ���`TdfR��,D@�g,�����ƥ@��3g�����!���[b�z7U(�ql�Z�/�`t&'
������y�8�e'b��&��}��д+���Hc�Ej�	�G�/�Z�o�.�2��8������ _jZ�
�q�s�-�����������=4��Xb�e\�4Gfu�l��N53Yp���y8�	*�5v7�e�z`�����f�W��J���Gz�!�{�/�"��H:I����D'|o���BSr_#%˺��=�	�\D��5�����,�Z�����K}@��/��-��ȩ�����X���6o�s�4'z�i��m�W.��]��Tȏp������L���ypb�:�k<�rZ|fz�u�=���w�7�I�	�����
����D�v��>���͗�,ɓre��+IO�|�I�0y��}�x�m����dz3f>C�u�j�~�V�E(Y������ˋ�x��>�|/�)��_�1�+�y�-���)o��#ߡ�bV�k��'NQ$X8U�V2����;���Pn~���N&Yu��	�%�򗈛4"���`�>�x_�#��+��#}��&��O��ң��.*؏��׌