XlxV38EB    266c     90b?�p�����8��,v�䚩��4*�%"�X��!��N�G_��)��=Հ�(I��	��,HڟG׭V��~������h�J�Gp��R� �$����bk}�N�k�W�~�ݲ;��Kd�è�rN����(Ͻ�w���[3�s�4bS�#~��6��7�z�6,��;���q������ �/f�O���PT6�G�v3����ٞ�x�Т���:v�\?7��<�f�@�CՑ���ȋ	saF=�����\ѽ�<��i٦�s��)'�ȿR�m�p��B����O�=�K_8f�	�����)����[��k}~ /�0��t) 4�� ^z`~���A�2(M5�}�;��<͇�y���/G{e��fl�N����վ�ĹK��V�G����s=�W�����=��]mxf7�]&^#?����ꬹiҜ�����~�2Gڊ4�Ͻ��e�%��0��ׄ�F# ����Cx#�Y��9��XO��'q2�������=Þ�����&���U�ˊ�G5����T:�e��,D��DsD,�4�?,bP�K<#�:��sވ�D���7X�߰᤾__�&:	h.���f��v�C����9��@�;�!�Β
�����zK��*���D���_k<G���*��ǳ	$����Gگ�""���P�n#��Q�0u�Rup�o>�;��a��H)�(���?<�®|IB��i�E�����.w�J�_QN�[����!h�y���<G�"�Jk2	���w�b��}�8|NÒ.$�w�������������,���K��Me�����l
�IEN (�Bx����0����2��Xc�VM�*�gq�o���U����0�z��ـFq9F�2���R��ʅ5׮S��B�m�+���y�.V#�PS�r�RZ_���k��F��Mw��R�X�����=�yf��'��6��l�=��4�x1\{B�D�S���k3�wW��b8�߳XJ5�N:�UR����	��Z�7�T���ʳ�j�iX��)��ь�? ��.�V��d��.��,�t��ر%^ƏE"��z�=�L܂P�␠���P8�o%�	?t��Ұ�X��)��������-��Ep����j^cql@I����˰������uc<Y�V�1'=X�PI�	�I��7�{���+"�zF�!K@%O@����&J��g����� �\Kﮔe������k��Y1�g�^�R�����[�eH;��F���o�O�xqLfu�)\��5�ѡ��&��PQ�aEy2�'����M�#$U�,����=�$�ua&׼���ā��$�.��A���������2��k��������`�Q��L�@J���	��b@���b.f�&����
��_+|��MH ������1LM�m��?b>5�@��`v��榄�����1C4�����s�n�ґA/�>{���G���p���f��JOqx�g������me���C�j�Z^��f�{�	pN#��]�-�_� @E���ڦ�L9 "�R\I�}L�Uo�Q:�$_L�ѱMxj})�]�f�E���6���Jm��8��\�ݳ{�����_h�Ék��t� ^Ѥ��R]Q��4��h��nd�J�R�5o�`�l�`+S,�����}�8:��Ɨ�Ė��sD^(������%�v��с'���3�����_a�T:_�Yߥ2ZK��7� �B�B���׿{$u+y��Q�����؍ʵ�Y�Pp���+�^��>b��`C�v�$"+ǽ5�c!%�o
��qd9
�(���s�����~�(��G�\����k	j�a@rKV����Q�z�L��Y�0�{BӮ�"�_�KA���"��*�w���3ϺC�����{+F֟���l�R����u�l�Tv�_�}g��&����3�0_`�m��.� ����#�^�<fS�$Qr6Ҽ�	������8��^�'Ϩ��6���E��z	�V�\>���T[�sM�D�vI�t)�����+����2���cme�)�� '�c���s�I(�^.7�Pޚ�
{<c�	P~�-�}* ���
8�5�o��k�ۢ�@@��n�`&��$�M4qkcN��s,��tsF��GI�����6���y&n;��S����QK1}���C:`2y�3@&����}]�� ��Y�@���\!��&�8/�*�6I���r<�Dc��i��oc	�[���.��㳨W�^M5��m�: ���b�6����Y�It�,�������U�Qi�