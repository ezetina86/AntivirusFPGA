XlxV38EB    126c     4af�6j�-{`%�P6 �8#�����UZ���$����gU�S���5�m�:a6��l�|}Ìh;���Kā�;�� ot:+X���?��ƒ��@����z-o�+���D^*F�k�-���T� i��8��Qć��T)�z[�B���s��dS��>�غ'��ٕ|�cԔ��++�1W��v�H� ��N��yΗ_�L�)	�Pv��Re^h�N7pN/?�����}�V�(s��h���O���=�R�[���A�`��� �ԡ�>E�P���.���fHV�|�/PD�HtAE5�z�!��O�S�v��qp��,=�+J9�w�3��%���+���ȼ7���/;"(%�)���H��b{:B!~F*k+
�L_ɫ0>�_����N&ca*W�x i�}�!k(ׄ�RM�[���S�����GzQE����h�)|�u_#��;�����|Ng�`ߴ�F�l�\-��)�c��(i8z.`�*��5�* b�f��:@𬵥�o.b��C�<��&9$�>�0��� L%EL��uD��7��;kZ>����c?��@����`k��t��@؂�O�L���ɍ�8�����O{�B�Ge��ܠ���������+ruzgN{��9'�"��t��<$��ZD�>.�֜ 1� ����N��J���X<�r�� ����oAv�R"F�;�W�Ϧyd-y��K����B�U)�>o�y>��YϪf҇c�՟F�R�l^)|l!pXf�	�QC�5�����t����.�M�N3�mT뱰�%1�0I�G�㗂V��qU����Z�������Cʥ�?�dSL��i����:L������ȱ����͓�����Ul|�� ��Hu�s!um'v����ʲ�0�[I���V�_T4��n,�zf�1�{��y�Κ[�w��'�؛W&��M���/b��8�$K�M�i��c�Ͻ-[�LMC�&� ���{;�Z��A����宊����W^Ÿ'�L+�����Xer�-�YOd��ĺ��>�ة��Co�,Dps� r�"���yQ]1M_
�	흕A����r��dqP'�����%���ېA|�ns{SÕ�D���$͆��/oΚs��֏,��+Quչ]@���^�,\'8d���/�A��-{�������67�AsC+C�(p�<2O��^�� �gU�