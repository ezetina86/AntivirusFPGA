XlxV38EB    992b    15e1�$���(�,�� ֆr�x�TDǜs��O�)I�5!�b���������5�M��p�K�#�!^�j2Q�"o�K��9[2S���]���շ���^��q��~,S�@7\�3�2���,��i����n�dC	/k#9),h�=�����R�{���?���`
 F��{T_��_c��w$^�Z�ltb[Re���8+�N����f��J5����^~|�W�]G-I�����%�O��%��2�;���t�՟!M�f�i��B��鯡�?hҺkA?U��2��s�΂R��\�gr���I2M�����5�M�T�����a�p�^��
5 �o�S�Uc����0�\�� ��&]sT>)����Cvb�{���%Gʅ�����F������d�W�m��BĊ�[NH�c�)S\���b�}E�Ը�#(��{�'4���ltw���=wt�$�g�&��mif_{����gvq>n�	_3ǋ�/�b�݇�]���Sf���v�s2k���oc��ȱkљkƺD{��lE<�ySͤٿ:NF
\�[�c(�<�x�(�[��F���$#Z��}�u�0Q=G���������c���5����cu�ywh����`�&A�hR1���dL��3n��~�A�L����C�6s;.6|�&�|�
[�^Nt!Z�k�G��Qm���j�5����,��r:�DOH��;���\{ٌ����	����i��Z_����$��Z���N��¥��n���������{��5G�;̵�H[���N_�V|m���j��|ݦ���m[�D"�kn���t�dKL��C8M�W����fB�+���LY>�)c!Y"��z�1��(���D~ ����73�&aԫ<6�������&�GXۇR�mV E�<fu@�� �G �lSɿ���u�o�0�䇵L�y���|��1D�WgY}��,-'d�:o�
�8� ��שB/�
����z�`�:=y����o�Nz`��������QH�#�#]���lC���g�7��#�8l����M���'޲6�J�@��R������Z��
,��"&4`"ܙ�/�x�A��=}���4���T�Y����X������i'��c@ļIF�%zE1s9橉D䁤�~>�����MV��txI�03�~y�\n�7��	OK�>�c��"p�Ḥi� {-@�O����^�֓����C�v��`m��ʲH��VL� I�x��@����ҡJ�,�"8(�׾Iu��
i^2�\���f����OG�2��v&��~.B���6���%���ݷg�뉝'��������[ou׫����=>���]�^���)`s8�+�B�6�z�'l
�����;_u����E��F++X���l8�2֛u�ӕ	ь�x���{��\��md�%։Z�u�p+L�:����(��Ht�eU����;�㫀�{I�]����M������S^OjƺaG&v~���M��'R��ww�t[�;Y��J�#/�K���v���ص��6�oo�}�V���-�DH5kJ�Va���1�'��ce�g��:�)��1��&�e�)��zo������7.����G%�������v߻�/u���n�_<��)����3d'��0Azn��/3ٯ{lF�#ET[�W�����1+�Ȍ�@��Ue��o�rO�9��N�y*�b�u룻�	�Fr�W�f�ۜE�Y��� $Qb��K�u�oē�V)$�Q�۟?�m��0t�+�߰��x;���fv{�ȣ1�¬X+�7�\�����Яo����]��3�.ufZ�u{�(o�Ȱ���bކ���y����V�l3w�5��x���[�՜]v̓!�V�%f�c�FM!�s<h�
eER�~YӠ�� ��uټ���]���E��ci
2�Y�o��H�9>����jc���y�f:Vj
%�TCI�1$m�J�� 	DW������4��B�[˂"��#f@�L���J����s�^���G�?R���K$�n�/�:oJ�c���'� ύ���Ǚ���Ɗ�}f��ys�����+Z�B��Gn����gK�����O%R�y�;cQj���Lj��"��
�l��>�A��t�>�c��z�I�ژ�םL�)1���j}Q>F��Ĩ>m��?۶F�Bi�a�Ex2Mi�)���{;$�>�āy>���� [��dgzI�S+~�Phk<Q0L��v�DK�� ]��,bv*�bƐ�m�f�cj�E��ݖ�'Cq�W�F�l'aT�f+P�5l�B(�mS�H������#�|���OE1`��ކ�:Va?`.{G�b
�#-;�
T ��\F��ۓ-@=gJ��+�2�B�F��-��1�@�i7kp��E��T���G�[�-u�7:N~��Y�h�=2��!U�i�x?��S�
p���1�.��������BSDZ5K}9J2��j�l3ɝ�����T6�+�$�n���t�y��M�Q8w�[�6{>�E�v�r�����pFMwYTN�>P�!��hv�P[鷔�[�����qRKB|�����t���9qP:6�����_ְK���!t�r��߸2.�+�v�N�DK�)p;4�V�hp�ӣ謁B&%{�Z�^��?�? �&W�դq;M���	◤-��������w��-q���#�1�/�Z���A\��%�����2���|�n�+���h±�F.��lȲ��z���y j��d�¹w!�{�I��bFJ���ضR��Zm���*}��pK� ����:�[W�.��[�6�:��X��w����I�0�ܜϩ�L�?1�rYI�Z������S�5�[d����e@���������8PgxZǥ���θ�{�}O��ो�|V,[%� ���*-h�{Yn�ν$m襁�jK4Na���li�KN��KLH�/�Q�.zY�l7�.҄=�jN<������|+����ac�����Hi��r��m�ʀm�J9�=o Z�]�S�E��N�=Ӽ��>y�V�|$���t�g�U�
�F��Ʃ��:Bv)M���bʦ�� ���*��$�w��n���ҽ%Is��@���t�|,g�g�מK$0�Oݸ����)�	����=rM�����������)?D;	����w�S�BǍ݉�v��$�K�=R��o�A�<n���ᠿY�AՃ!�xH(�Ҭ���,�mr�jz�xǑ���Q�\d]�A��Ȟr��r4�#����`�w9��������F �Fa�?}TF��O緙r%:~��8bt{���%kOV:�P!q��S|�R�Lz��"l��#8Ri$��Ev�]6��*�P�ݥU�	�ٌ�-~ɡ�c�!0S1�un�+���o?��MnK󨱈)�
�f�h\�Wp5L"�[ڈ������v���t;R/�V��F�1����3��p�@�	�t5f�=	�XX����->�)Xl=RR��啵9���ZƜ,R /��i|����=�d�� ���X9j���i8u?g�W���4}�����[E��b�6GM��8�$-ɷ��UMg���`�?d��M#FA�i �)���Q6�������HIK��L�R��M���󩯲&��4�5K�1����u�ގ�V	�`�h�O�f!�;(��53vv�j�n�A~vfdSF�G<rBο�ɝk�h�}iB�	�9�-l����Sn8ǚP"��/1��^+��bW9�IV�I8$�x(�4��M�$���Ӝ��ڳu4���C6�aY����O����!?U8�����z���"W�ݙ���yv��>nm��"��7��wA=~1�u[�se�b�p]�*2�����:\`��"��`�TIA�0��2��xϚs?�;�Ze�E��mD�&l�n?� ��ޛ�5-��#�F�>�yy�FŻ�'1��Q
�P,26�x$�P���d��z�V�k
8���]�-� ����? �w�E�g4�Ƨ�P�n�G��OPq��HS����_���b%~|*�V�T#���Ƅ��N���0����Wr�M����f%���pR�>��T	EA�<=(�@��N�0��ę���b��S^F�1~�H��	�K}�x���dBv�����}<�CX3T<m���S 2�(DTţ��t��i��UGX���x[um�?���rn��Wj�pu��aC�P?�ur��W��S�sEvh����X1��`JB��u��s�d؞ae�U���Qr뻽��ՠĦcֳ8�o�#F	7oz��o|���!�}�m���ף��u 6�+��ֱ���'�;gw�F�g�,�7�s(�P-��<����z�.7�vd9��2Gz3��6aR� �+��*}҃����4I�P=����Zz��g����Q��!��e�g�Z͟x} eVj)�������ƽ�-�'y�a�3#|�8NF)$چ��5�\�`�.���(V4�e!o��Z�1��Ώ�qO5dݚ�m+�С�896̡JWR��K7u.���%�<`��\<�Kv��O�V��;�9L|m�1F*]t@Ю���UW���)�^v '�/'���R��i��D��hjm��'"s��6�N��J��liy��)ل�\כ@�Yp1HV3[G��u���#*�
Q�fz�|d�,g���[Fn~?�`�^\vj���W��|rc��u
��-��ɵJ����jw�4�7Y@F�/��J��B�.�[�ǯ���rO?��N%:B���)T@#���V/���r��p�2]�5;K�;������iN5a�K�qK&_m�؎:���W���U���fR|��N�ۋŌ�F�"Ne\gܐ5N�xΣ��� e��r�I����xWدx��{�/�W"�e��Z��S���5:0����̧�3��c��q��S�M�:]����ɉ�=#��V&�����[�h-���
��D|D�1�fv_O=�R�Z��E�� �/̨�ՠ>/鰙PO;1y��~}��Um3~��2S�8$�V8s�`��{�a���	A��E+a�}����g��-)z�T��w�dv�����f����JC�B~ߏ�1��"�v�����=��^{����R�s��U)t��=(�"�����8`n��B��;|��h���E���'`@�?g_�J����F��(�a3���@iV�1�i�F&��K�\��Z�r�a����S~��ĕ��#x[�F����*�i$����ҟ�X�{N���x�j�\�P��[IǴ�Vk�3ʅa�4V"1A;B�uG5E�r�+�-�}[57Jf�^�?�Ÿ;_8ͪ6��Z�L�Q3nO�GrSmAjM�ܻo���?QjR��9��Z+�҄dxH*�?X6�_%Aq�s}�aU���-�5�B�̮�#���y��K$\�
�:��M48Sw2�h��e+�j����k|��8���Z%�$�dƘ"�������/"���9Sn_?_����ePWvV���.,Q�^���-�S��u8k���z���2���b�_Ě�#R *#�Vw���<�(� �