XlxV38EB    1161     48et����|�l�H�^ޤ����u��w�f����qF���2��2G��C1�Y<�Y�uFw���)[?�)�A֪������#�loY�߁�s�¿��d�B��֯�n��d'ғE�ޠ��m��ӯ�����V�����(ޛ���t�SjPOD�Du���Y̑Z����i�;,��IyR�~�pA�6wU+��ax�8��Sn�DQ�4T��	_��n.jH��#3/�WQ!���/��q���� ]B��<.�y�U�d�%��O4�q�vgA%�~Q���bn/r�� Q��\s����Ϛa���XQ �e=g��ϲs��REh!�b����N�zv7��}���	g�i9�҆*e���|���6���X-�GU����}�[Q/�sZ܀껳X_�6����+�|�?�	��`{�"��+��-�!?�=��:p�3�����n�B�d�Ҙ�n�ZUH��yB���B��ro�'z���pW�耘f�X��%1�$b��]���� |��&O�׿(��m�*e�!�نIϑV㾹� Ъb^�[F-�Š��=����;N����kD�n%=�ɷ0#�ə��#�q}��q��MQ��n���@O���~��:���������l1���t��3���	V,|&6~*�cT�h�i�	U̶�3}��=/U�#a�*��}f��X�����)ȿp�1����\���N�
��^6d���^�.�􊨁w�u�tc~C}>�Tף-f�Q�bQP��oІؘ��WC���ar���1%�鈆���jGGm��μ�~[<SGx��=���c��{򝁺w��7謯�ԝ��'�S�"���CKP��Ξpt���c�2}�`��<U�<`j&�@� 2 �E5��:}byk��<59_���&[k�Z���1�)�W����xL_F�,��ђ�rǂ"/C��7!f�����J�K�F*��"�N�Kٸɩ����@;K!���I<��.3�M>	�E8�ƪnw� �uDs��X���I�HG�\��g�>��u������1c�t�So7_��&��������A��)j5�W��������z��8�/!�����#5�������Z�0`�Q�)��t:�K�Ur� |O�?߾*