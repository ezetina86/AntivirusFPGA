XlxV38EB    1def     551v�4�`Qu�7�_�K�T���mjN���j�#�#����N�-Q�X9��X֡�}X�V_����?�5MN��u�K�<E��3��fU�ϗ�cj ����H���ƕON7?j��2���W�����\���ұ���q�w��0�]�M�T7�m�?��{#l���A���LO$wV���l��o#\9�>Vj�XL,�ne��P���k�V���L2T����vU���ͺÛJ�h�y:��+C#�X�*����v�;�������&so�G^��~��p_�E�ujM���v�rc���2��x.�q�B�x⁗�f1�z��8/b gb��O������Ɠ�z�p��D��镈Q��n��-?��cg����t}F2���Xފ�@y�^ ��N�>��٘F�TY���K�͟�wZ�jU�8��ҕ/��E��_n)�n*gsrJ�أ�hh/��?h�X"�y?ߏ\i= �9��r%L��M���P�t��I>�\Y�f���>�V�o�c25�b����x
<.1ΆzN6t��&U�x�]��r5TX���树��d?����9"@�If��LÃ�x�F1��o�ϼ��O�GH1���Ok�zQM渙�Ы����h<���ȯ����� �	�	r@WQ�/��l;��l� �֫�Â ��C��Aƪ��W M:���b�t�-5��`��� �6lǬ`�ʄ�9X�Q��	�C#�g�b��D���6��/|�Pt.2
��-�u)�����
4��r�n���į_k5��#�Q3�N��d��/��N�)w�;��͐`��^��<�RnP���1O6��N�z6[\�?P���>�0��4��P�c�G"u�����0W:��#�-�u�-O�l�K�T�~5�SvX¤��(������KX���F!��R�L!E��.�}/��;�<��X6�v*.=W�5A��_$�m���jc�o�0v�+�1R�`�����T����l�����O��,�.FrǛ(kqP4a*s���8�A���P�vU׮z�3�|w����������/Qd�x���1�p3�A�l�k�� %(����ȿe��H�.�D��r<=VcQ@z����g�#B[�x>�f�����0dc)ac�6�0/�5O��1iD:G��x��V�	�fh����B�+���N)� �*x�wv����7g[���yX�R΁vz>U�܂]/U�x*�/^�G�sBT�J7�U�=L��*/��G=��=U4�b���7�{��f�fj���-Z���&!t�i��~.������e�a�T��*���j ��c�ٷ������˿ PAz��