XlxV38EB    4ef4    1115���4"�?ޘ�%hK�:�1�*^���-��O@D:,�S-e�ުL�w���rƎ�]�?z��?�e��ӵW����j�7���a}��ʓ8�y�f�5���w�._��T�.�}m��c��2�`9��q��6K�0�#���7�����^��]�-��K&���d���RJ�{�)^����P<'�+y�-� V8���.r�di�bUf�����<���
ծ,�,�3�d��	��RT+����ʉ�4���V�c�sاHX��4����1K�7k��<��'D !�N�>�f���Sl$�P�>��]A����<x�P(-��X�p�qQ�����sM�2,���A��?ۂ6�߱�C�`L�f��K�e}c��a�νV���P���� ��}�S`$�`]:p�&���,"D��?�k��l(�`W4O������L��x�u%4��@H2;W���۶Ӡ�~R��y�L�҉�zd�BZי��D(�(ӽnϤݦ{Ooh_��A� n����)�.��1�7O{�ze�}F�k��bܘ��t�_�\!�s�JhE�~�;�S�p��]�Ԏ���4��gؙ�����bZLXV�5�H��쌮�ƌ'T�7��J�^$�'P{Zx%!�N�|ј�i��RQ���=�Sio�K'�|���4y)IϯњO	�;�6� c���rc��x����(���6*���U@(O,�����U_�
�ᗈ�9=�D����3��D%k�����y��=�<��m�Fd�y���6ltW���+���1�� 2��*\�=7]X�=��J��v8�U���"�� �&B�C��#�Mģ���z'�8yw*j0y���btSBTۢ�uL��Ql]��������5]��3hH�� Q�u�!��9[�O7���b�rwR�f�ES�a7��'pP�e���G?����L� �[z�7�:��ɳvNR�Q��x��m�=�]�愄,���n�=�Ug�d�������8��g������m��ǾkJ�'3�8�]�ZmȐGl �I"�z���mc��+�d3���`	��#H�a>��\��R�#_���|��euSܻ�)fd�ӗo��y�@n���:M�e��q�m��,��J�1BK'��dv�Q驆8�����v�VMVkt:@T[-Piī,��=A��Ԥ4�(����D��{У�O�f8o�?V�k��8b����ɔ�ў?�<#�vT�ɛ�/��w�.���k{������"�ҵf7������X��y�O�׺2�޳|)9"Oo��֞�j�Y�c�{���(;��j �<%?������sPY�>>.ӯyc�/v�_;c������Kb����HjL���]� 4��5z	�ZA�d�.D�d�kш>¹�KD�)pʩDu,"�&���s@�%i�rj�*B-��[��?(���z����
��Ze���qT��l:6�٧�p���#��ɯ��/�Sϝ?D�ŬwGн���/�s���|(%�8$@��Rv�R�25�[���>�C`����%�o"�+L[�����O�j�k��M'x����u������Gߠ����<V���t'��R�G��OR��a�OPhT��l���S){�d�-��S<�㟶aM=v�-���k�"Eh�_�Vh��Q`>QY!A$�(�u�0Aa���8�ê1��քt�'���5%-� �A�;�j�өv¤mzJ�vH��9s��W���z^���!�Uu��LW�vb�>�y�N��i��C��!m��.�r�P�u�f8G��6��K+�(#�Iy��#�F;A��C�`����ǻ����vJ�r%�[�K����=�n����>=MF�L���	A:�KM�}p�����rE@����H�H8|�f�&'�~�����--�!����e��7#y$�����~�I�X�}$Z��	)�l��I1�K��!�� "6 Z������	�uo�Kѭ�w,�tH"�APn�[)ip�53�|=V���'��^R.�g�Oi����\5�~��L;�Ҷ�M�R/�QG�K��]�=�(\U;����l��W��}
�[]��p2\'ڹwT�eErm���FG�a����ζ��q�`K��
�A�㧺a��1���s�j�:}Oi�߻���P6A�|܂��Zi��%@�7z�eZ�^\�r�g'y ���z�ߖ��$��hԮ�rK�$`w;OƓ�خ�;�p!x@�1�4&���*�u� �%��nܞ�5J2)�WB}l�6�LHԍ�75Ǫ��ߊ����$�^�0P�f�YE:���4����3�b���F9{�&g|�8����?��y�k���֐�fz����ʥhbY��(�H$�����𝯝�o�;E�ke�a^�¯�)Dc����p'�dp&�~
���
�u�φ��`Lÿ�c�˳qY�F9��W��5B�\��*���������֞\���EU���RS3)��GS��,�@�o>���8�����)*3D�JY\7�^��5g%�-�B�p�#�U��Œ�)�u䢟*�����7Ekl�i��↹�o-�4��9�J�(%2+#}0	���w�ʈ�?��ԁ �&j��eWh5+ࣦ�A��I 8]�4$���:��HI9�nIW�*��)�-_�Y�	���S�Q���#U���8emB�zxِ ��V5���;��?��n)٦��D�	wV��}����W�1����[#C E'U��c^;�(`,�^��[o�L��n�P�*fIh����(��wd����L��%ب �<��MA�׃�/T⻖sb�B2�,>r��BFjdfp��>�(�΀��H���9��OH�QsRn���&��t�$��:UG�p���`5����HƊ��r޵Uϫ�A�@�mL:>$���������	��V4��@���
;t!�D�wF'L���s�GRb�o�BŃ��p{�3�'��R��v�������z]�
���^���:��-�H�^�㡝^!*ri��i���z*�c�Ŕۉ~�q��G�f���)�))`�ΞM3�� UFMd��e�Zt�M�摑y��S
�չ]���t���,�����F"XcP��X�̿��cx}~��jH�-�W��rN ^���q�10�(���v�.d!��>�.$��-&�u֧+�n΋:]@����=��=#jb��iV���{}���>liܪ��D�b>�6�A�����.�i�:�o���J~���3������B��S����7NLl9O�N���U#hs�2:���M�iJ�8����1BW#��l�}�`�1�EV�Ͽ��'=Z�js~=�F� =c�i6Y�ۖ� ;�w����s�r=�C	bmX��Ԋ�����;��x^O~8�)�B�^ױ����*8|%4���hC@S��j�e��_�����s�~�onb�].!�i\�+D���*6"^`�7���L��9ӄ5k4�Nc�$���a+lɕ������|>o5��Pp�DP�db	�z�*V��K�aWV��t�#R��]=
�G�;���P@	
Y`��v��< �h�Dr���K�[��H�NaY���<[���M�{J���|��hC޻_��o��
c����5�nL�OӨ=��V�;u�����o��`� J�[{�./�o�J����潦-�\@-"g�\F1�-�]�V��Go��7#��%����`=���y۸�!>���6�o�G� Q,:֥?�|V5�X���bs5���63=~�&��H̐��iZCgL��U�sm\���?��=��)��s6�M�
۽��O1uz�pS��6�4�>��+7�4�ʷ����W'P2,X��q�a��emd�[��fӪi����p�;:�1My��i��S��s^�m��dk���fCe�7�҄F�^��sLV�bk�K�C ~�,//�;��O1m��ҽ�����J�����6�z����IK����	���K; ȕ�����M�.���j�~7�K�'�(�Oylsw���.�$�l*�b�TR8[�~�]A.]E���/Z5�T����0B#�ء��v�����H�L|]J[�'���%���p�-k��/��&���a�gb���$�S�=x�:HE7���u�_{��`����Hb�1��N`M��R� >h����Vpc�{YF�����t��'��\0��s/�a��f�+��_��4)u��YH������Ol��h�ߴ���W@��n�Q9�pT bH`��IxL���d��;�'_~B9"t"^�����B���,rݪXny_������6uO���h������Kشf'Ԩm�Ze(���)Z�;6��