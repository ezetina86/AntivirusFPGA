XlxV38EB    1168     48c�����2�7%�=��ٷ�5PI8���?�@|��Sy�@.�������m����M��e��-~Z�M�%����Ш�	�h��Q��e�/~�����i�D�$��a�m����t�`�O��lD��IQ8���[�>�`�(�`����>9:h���ä2_(|�/,h2�3#�S7R����N٘���z{鞄=���n������g��{`Ť�Tt���!�%�OCjt�X��U/p)�.����\*����R2�ߤAw�Dƅ��2%o����.m�w$o�>��e	��)�^k�͐��w4��G����<����1����� �FyP$�:�"���hc�[1���oB��2�3P�v��SW��q�A���fW)D�C)I@����S�EV��t��"b���񜅚:��q���%W��1��P;����b����<j�<y�Ia�;�)I+#W�l������S��X3� �%�|SM�Z�����[֍���Ɗ��.>#5.���v<B�j㿂%`e��q�FR�0I#zf����U�;u�h[*�3<;���N������!�Zy�t�N���1�XA���4n�\�I�-�+N�<U*�gW.Cලރ��*m�P=� �V%4C0��}��Rƽ� �7Ђ&��ˀ����yڧDsث�k�k�.Ӌ��_����䳄�4��4� &�;�#J���0�0�؈`�E�Wh�"�TT��>�����Q�SQM㘣�Y>3S¦���o��8���h1�T���|��U���Ԫ*~�=e�Ra�u�Ds:��F�+&���)*�v�P�3y�)��#���y:���E/~z��"������ϒAHU.&�>B��0�v;�6��Ђi�@e��_X�4��j�5���j.م�<��Zy���,)NԱ$Q�������]Ei�qZ�O����qG��S��z��T�͜��w-�ڒ�٤��fu��J�j�a��xx�;�ݎ�/ga2�yt�D�uT���i\��0��WpD��D�E�v'�s�O��ִZ��^�>>,�t%N���W���'���E�-~�S<]s�U̜DZ�UB;�� ʣ����,P�V����vu�`1�2m?��CQU����L��9b�D>�ĩ�$|��Z��<-p