XlxV38EB    4aa7     c33�o���1�Ef�Q
d�u����=�c�Pp����]�+"0f�a=�T;�L�-�Z�h���vua��X�!�R�JA��N��H'_-��1=��_�GWK<��&?n�H@���0R��:i臆������T�bؑ�9�.%<n��3���w�,-�q�p�cʵ�+���z�}��;7��u�0�G~��&hfv(*��{X�,Ŧ�r���W�9
PNP4 �u�%�0���p����/㧂��h�T�4�0ĝ�{�犳������_K�X1�l���m��eO9f����R�1���R�mzW#qQ��B���������t��z�p[��ɴ?\�r��O��hO;\��>��|[Y�5����n
f��8�p7.!�B�&0KC��(s����0(���a[~�������-�&'���d��E}�ր�o���؈�UMH+8��;�sC��{�"Ѹx�Z�_D��t�>
o��
�4�'�3$��hAb���T|ʾB
_��X)�|S�ʖ�n'��y(^uz~m�i���)�@����a��<�͵�K�o�=�%Z�V�����iM�>�ٔI󟴡���"b�~�5ۇ�5�h��SK���}��HMݨ�Q��z\8�+��{m�Iw�@�̑��6wc�+ou���F�w
��+GJι�f�X�]NA9�
���"1���{���b�=��6_�u��Z�B���(;MT�KW �����Ɣ?sw�����ඩZY�F�&62�j>wB�[�:��Vʊ��eF����sϜ5��V�D7\��
�W
`wr�����Ff�F�o�mg�#��*���Ғ�e��m��9��\T�$BOs�{T��%"�i���Ҭt#�����6;*əK�=O� �R��Q��\���U�}j\_���p#ԡ��� ��Om�I��m[k���� ����|E�;�U�	l�O�F�9UR(��e~ �-֩�ƏO�$��ք�q�Yf��xEO�8w���U�S�B�V�a?��h���S�O�<��|>M��\R��6�!MϠ��=�q��;YCn/ۨ��
S�W�ƿ����[���-q�(��� y���Q ��-��)�_�ܗ�cJ3�����j�ܞ�$1`Jк!�Z/J�7V�=h��&f K"
������YO��w��Nay\���9���<����rq���L�E.G�G��m�Y�i���Y�a���<���^� vH+I�
39�
�T+�����q䪦{D�u�ې��ʱ�fo��e���|��p�t��iZ~�i�����$jM�1`�^�E�u� ���3\�J��i�
B�g��W�=3�U�2Pm����!q�C��V�4�+���
���H�O�h�;�M\#�P�2�6-���hs�zjb�ے�p����X��㣔r�H��^3�g�ͽS��t�$�:L��J���Tβ�㈝�w՗y9�a�a<���f��s~U���ܥ���?[�su}��4�S����$		5�n𿄮�
�Gkn@��ֵs>���˗�`�$vz
��zS=Ε{Ύp#$+�W��+��A����zU2�*��c<���mv��`sX�e:�����hh�I�NZ�6��Y�ڹ��|/�ۿП�Db>�J\��>z~�VɅR����QD��^��I��t����P�9��F4��}L!�I}�:�yr�O!`8��YL[Ɓ���2u�G:f���� ���P�(AP���i&*����}�C�s�t�kk7�Sď�x��lu4VE�/4���/�8��ý΄�
����^@L!�x)�_���n=$�;����z�B��C��"�����6C\V�P�nN*[D<};5�{T�Wa{j��f�xܠ!�i1~��[��F)�����*�xk�i�M��L�O�߅Fpz71gꝞ�B%"�%ud�����VTbd�*���{�z�TBh"A>��h��$�I�H���(�`���h���>מ
�B�G��i�2��"~�3�*]Ų�>�j����!�o6Qb��W������G���75�n]��B��h�
e�ILzg����r"(ܟ��c q�j����vs٠&ڤ��3"�����S�W+�³��ɏv���;�3 �!SNWI��O���l��R}/��
���@���ߠ_#}o��i��Sº�i����>��.�>�`���WY�J����M��J$�S�ɮL�T�)k���:�c��m9�.�����k͒8���� K�,�Ĥ���2��o�J�q�zs=8}�)Ӹ!�>V�����O����m.X����w�S*H���T�%���S��Nk�S�cq8�����f�e�����zK<��2:��������x)Ɋ�@ ��J�+�*�r���c������Q��j䙽�K�V�3\�h2���P� �p�ZUnE�|q��my%���y��������>���豥[֭�N>XebFJ9�k�X����	�g��4�j1��񎅐��I�9��O�v�T�Z,�m����u�%\�T2�Ԭ�\ds"}��|���6@��I�xEV���2�а �����Q$h���a��9�Ĕdu қk�k� ����"���4�C*s�|vbD2�+��n��
���d�[�%;�K�Vs rSRq�.v�Ӓ��y/��r���̈́�i�16��{�uʀ�T�]wSX�JJ�x����,���?j�(�_�����Ɔ�e��H�y�u�:AH���D�ʇþ�����n������i��
��
m�;���ED�<iC"��wwJ댞�(r7Q���*!�i����3<J��Sn�.R�{x���;̩m��n\���4�kl��|Y��ΠKkyka��c��Z(�-W8���ޝ�%������d���9�N��-ω!���C	O�d� �`�"ڐNf���;�"NQ`*������՜팥������W�Pg��C�����l�@�z���"G����j&�GF���q�tUծ�X�FR9_����e���-j;ԧAv�UD��)&�����Ì�-��19P�;Ȗ�z���+��"��v