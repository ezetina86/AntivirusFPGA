XlxV38EB    1cb7     5e2�S��~�ُF?hpZx(�%V�?E�½1��
�w ��.�F��V|H��1�f;χ`�ҹ�(n������o����T�g"��3�����ˋ#�7>2�~�6�	z�R��΄��%=�,���IԌp�n<�0��#X��Rݲ�C�K]@t��'/����e��n=9�j�g):��3���&qBy�~���r���n�L��W������X9�l��{�>����a��u����K��ϡV�T�G��J�9$l���{z[�x!gJ�x|K����7���H�!�r�1I���T\��yD��4�]db@4�G��=��V@�������7��z�HW����@�4ك٨�R�[�Q�=ޭ�����*��uk���j�ՕȬ�fg�B��{&# ��J9��/�Q���Sɮ�Ŋ�O9�J��椅Z�%����v��`��z��W&4��	$����-��T��b���ȖJ���N2:$���î/�~���DUS%�*�!2f��.`�_~Dܠ�;�S�&YHa:1����ڗ�^���.�O��WD0� 	�&���Ce�B3mNe�\���M7������{h����v{�X)��W^p��˄���A*7��K���`n饡��r]Wn L�^��a�~�/���,HX�ޖ�'R,>���'�� ?�2�M�q�q��3���I���F�&�r~��(��ڳ����5���0��[Z�o���_�z� ���=�T��"�@U���;X���-��ϛ��.他�$t~ �ꃳ��`�m���_;+���{��"҆_>Ʈ��<��+��9@�b��hB?��X� ��z�i~�?�y�z����`V,�)�=�՚ Z�:�ԨY�w���ʪ��{Տ��c;ٷ��r���a��Ār�?U�Ą�*���/''$��ƥ���rNƇfE����z��z���	��� x�b�n0�2'����-��K�w՝Mm���@j �������B�<)�����SGL }a���F�~N>I�Io[� Pi��*��B��z�'� �v"�]�8��ۊ۾���aZ'=�Zm qL�~HkC�菀{���G
�wM$�^�y����mM����/l�8����L|����_	�.���1�n+�Éf�}���ThC�j�!��2��<Dҏw�Ţ��W����`�v�(P�#��NC��:7$�ˇ�&�x���oX��7� ��[Ѕ�c.dT!�i�J���g��{>���%����uF�7c���lA�J�i�4�$�����ylaoR���j��'�y�E_��i�{��=)@��B�v��#��O%�V�W3V��#��������d��r� &=�h��3b�rڟq)��Ep�I>�ʁME�%F�s�|]��go�0�:wG����ղ�p��ƂA��Q�QYV�l�� �64R1x��t��PLY���G�bpjd�Y�ir�1ˍ�q5ǺrΦ܃.,B��l��P׵