XlxV38EB    12c4     4d5{�æ$���ڃ��a�_�ĕ�o�\��nI�m(]��b��[�#,�� r���0����t�7�{�?���?�T�|�2�����Tւ߰)Cgmyh�~�V8����͙�W�h��LQ�5�i̡C$��J�a�� ��o�ݻS�U~KQ����q;ľ�v����J�~����擛�>��#Q��y�F��y�N�2n]�[x*�&R��ޑ W�ד��E�Y��g��B�d�ةQ�5��m���B��H@KQ�Z����ц�.�v�X�?�k�%�ǧa��f2�u�d�v�4�\E����)2T��-��Ѝ��cAv�{�R��� 0�� ��|-��x��:��%��_�E9w�Ӛ��7 |tũ���s�,��M���z���ȶ�fBP}y_Oq��vi�?�P"�#�ϑ*݀9ܖ�JĆPwS���������Y\�?��r���j���ml�p<���D���#w��$��I��D)"|�t�=��BU`�l#!`�Ecוe��s��P�#K`�ٝNՙPظ�C���A��@Zo~�;ke�D�^�4fq��V	��f�OT��U�gcW_���da�� q
�>Gk$�@����K�ug�L5��]s���-�Q=RNGm���N*�:����҄J��z_RJ"��`3baą��f��OӦ���1R��[]���g��	ןw58��^)HTT��x���~���nM+���Gs���=�������\�T�����~\Cz� ����
m.�9!,:�a���ժ�~+���$�@��(0��9�:D]����,1X.B���kS%%��!��`E��_ӈ]b�~��Qؤ��UN�>B3 l�����;7e�Lo��;_���;��X�\�c�Khl��<� ��hI���5�M�D$;[��T� ���Վ_�����N��x�-�n}�@,���a��^�)�E�H��̖�c�R��~C�گ����0��m�M
�!����Ţ2A!5e��̀0���������B��ڐ��4�R@� ��yu�ң���z|�@z�Qq����+�Aüx�g���j�w���_R�ZK�i.���s�&�[��U`���i�~�?� ��E�m�J��}�n���EwjU���y?ઍ�?�s2u�Tս�XBB%YM*:��Z]e�/Z��S�%��RYX_)�N>˷ՈGj~�_����Ķ�}|�-"J���0:ړ+&-�-���t�