XlxV38EB    c9e4    1c68�����S{J��em�
&�����@D�$h)��˥
�,����w��M����\e�*��wl�UUQG2�7��U+9'8��IOd�14Qk�Q� ��a�F�;ƃ��^���5D����B�q���Y8�?��1�f3���W����[%4�CGQ�H1�󂍓DE�E�n���F%�!�*� �JL�'�y��j@���;�r͕����,�W���q��oNSSG�9|�k@���0ҽ���9�y���Bdv���ǘE�qtN^��rU:����Cm˳$���b�<���B�}-��['Uۨ������z����[Q^e>c��7���e�K���wg�(�U^w%�,����;��@K��Ȅ�}�u��x�{�����-ހ���B�:]���ߓ�9	oY�`�w�*��\��5=?b5DK%��~㊝�䘸�G��P8�m�a9KE<T��r�T�Vv��M��=E�k�Ĭf��|�Ɯ�3"�O7�mC���݂i�Z������<�P��rGݸ~�=%ЈY�ҧX&*�T����9�]Z�SY�B�G�t��
09O)D��n�;�lD(�/��x�<�m{ݏ��F#��=�4oC��G����5�mV�]�Jj��(�1(I�у�������Eݕ%��R��3FA�`^:��zG��v��`�s��.��E|G�޶kV�3���CB�*�xK�2�
��<���wr6R<d6�撿n��A���`���|6ܰ
,$��K�JLH�vZdu�FJ$���)N)�!eG̕ϓ`�
���3�ܟM���CM�Sh[�Z���ȏ��\�9<��jC�Iv
���C�k�&��U�|�����ۤc��I����:����D?�Rٱ`�t��g0�
�h;������P6�w��?{s�w�C+��@�/> ��2.1��6������WT���v�\ϕ1�ڰ���uƉL����e�}��+,���y�{²m�~�m��,�7���� 9yŒg�u6ɱ���긩Uq
�k'wF�&�]<��ſR"=w�us�p����l�����盬���{v=�!/��|����GH|rG[t�F�JKc��^�lc+@p��|u�K�W��|&읇�}����1?f��GYj��N����-_���Y�Q�Κ�=���n���{�_�j��Ȝ���c��c|H���A.B�����.�#��M ��ުޑ}�{E@��
���2����� ���Q�
�B-���OE~���㝪�D�����N֟J�7sK \j
�F�4��4����a�\��+�	h
1���\�y���s>���j�����~�8C1���佴׳�^�����e��p8�?^�[^v���0)t�h~�wg:EBJǅ��,K�#�1Y�X7�����K�u����۞PiK����1�{$
��7�4I���H�j ���`B/�=Ѻ�vJ�t��>l6�f�򯗖'B��@l�|�TUʳ��44���UrSb�.�1�l��%������-I��h~F>�y�3�d#�y�h{>Q��A��g`�`�	NQ��x~�( �a�.�c7�M���}so: c�A6�9G��T��=�~WCU֩9���E_̞�@j:�|kA�D��E����&MNcbDR�e�D`��zj��p��:\s���T�%y��	�f�FZ���ތ9i;x3T��Mvˌ�d}�H��{$G: �����)O�K���T��ӭb���vvn�>���J�O*j�=�����@���#��\�Y����?��=@J1i�e����r���4m�14�|#�>eZ#˞�N!u��L��jBC4vK��֙x3]W��KV��L|)�j�<�0R��B����נ�n�f�-�|����&�Q���2�x+,�
����|�9�*�?g��|��z�!d2��n��iؤ�d���]�Fn��`�w��b�n`��������kc{�HJ������9����-�uT<���[wN�RR�c���~����ζ�u*�q�J�]�Sǭ:4�/�Њk��gn����w�Ĵk��E7�F�e������ 5���~�1�ݽC�ɸWe�#���V�>�U��B1�<��6������u��?�}�)��k�Eެa��.���9C���231�F9��C��d]^���eͯ-��}��"ʯbw�1Vh�@y_��S#�
���?��-S���粶��R�S0z���ź<����������̾)� Q�s���(�P |h�i��$G�w��n
���>m�?��m�?�fY�v!���?ŷjN��Uj�Ҫ$�-Gc#��g�*ɲS*���r��1�v ��cY������q����b0}�Q�L�+$�U�lVy�	��3�8Nb#��K�+���l�O��߶�Q"�6N�g�=[� |��e��Pm�!�{I�,b�+J�p#"_\Zڔx��Y�V��-1�X�I{�C�q!Cau��俼����X=/�*�eyم/,����C5�&#�͉,>�!�T,�.c&qp jb��Y���bJ�$֐���!�
��ؗ�,��K�_��U��n�A�r|_/�7<��R���鬏a$��؜�),��u�t��I��%�%R�p1�9�cRfA-+݌Y�%=�ay�ue��B2Eˋ6Jʱ��<��"K�_��7��`�WH]գ\�P��'m�"�W���� +V�� �_�K�g�5a΃��2z8]�t�}��mLT��e�N�(�J��Tnv��`fE|b\�e%:<���EbB�����-=zi��h1j����N�����,\6&s챢�7����@q`�h�g�PPJ	�`ݗ��)n�a�V���jB��u��*D�?X���07����\�8%�O�02��ˊ&��ZՑ�b�R�� ����r�>Üc��([z��5%XI���d�06bH���q�c����e<��6g2����q��H���v�6?���Uk���}�E��C�6J0J<.|�����e$4�4{��]�M^�9J���3_���O�O��<�9�U$F��Y�$K��3����4���k;�&^���-��y\K']2�ө`���mo�w�'���|����/����wH$�y�FdA!Ճo�A��]6�v�j8��_��KY,;{�>����3[&>��3�8����@��5ZK����V	�$G��5��I��
\�"��H;��%��2yޥ���&�-�^P�Ď)݃�� �bO2�����OU�%4�pfK�2��.�k"�El���.��Ϙl���;�ͨ�[��z�X[�>���x�<̰͌�^��A��ާ��97��,����8�w����ջ&�y׼��;��WФ��ê�A�T�V�S����\�o��x\�j�J���ŀ��|-��`իe��E�2(�s �h���>���k!k��T(�G�X�|%=�Bܫ�>�bAB��%����|�R7Y8(�0yÓ�x"�\6A4ok�	�R�kC��3��K�G�3�5�5^+����=4�a�YxvXyT{A�&�;��D���?����U8��q7[`0�yxW����1IBACk=�h[!��-j�ʞ�6D
%sM)/��pQ�Fx�eO��Ֆ�9� ��ϷY.܊>2�0DaJa����gvP��R��/2�Όo�h'��*X�<�a�n�k��=DX����s��($v���}����r�x��/a!���������s�������K2_6�����O�X�Oky���~k�MB՝0v����m�8�~C2V��eŠ�%�4����ի���n���c���>�;4A��W�O��0PO�/�u/�����<=m��!G=�������7l����o̜�0�+�Wa��!
N���p\���"n�Ý�U��9�5�eq�W[\��s�H�վ��j���_ܚ�{/��ݨanM�69�Z4�G�C��E����[���6ۜ��쒴���6ٚfV�'S��e�Ub�L;o�@�n�C ��*	Ic��8�����f�P�/�I����]�lBAKQ~#�D�4fT���&��}0w�d�ɩ�V�g;u�e?Y
���5TrO/��F<x�o�z�5��g��8���]A�&m�@�l'���F�BS��d̚b^���
��3>MuK ?���ZX]#Z�.�?}���bL.�o�K��O�+���㴢�@%��Jc�=����rnc�D���B$03Zm�tv�^���x4��`R�N��m�".N�ӐV(0�>�^t��b�~�-�o�Ԯ]���x$?�]�z,��k�q4�[�%��Ypݣ\a�=H~{��Fn.Z�̀x4�L�;~r@�Q鲖�V��BV�^h	�5I����^�'�yڟ���s�V� ��D�a/��'5�[�>�#A�t!�g����x��"�s�H��ָ��!{N6��^%����?��������[J�� 5���^2�+�?���uF����+|�ԓs:�ճ�d���E�`��[s�R���k+���[?�d��h�}�fy_"�;�����t��0�_B�3�e.5�i��/�Y��V�Df5�=�!� b^i^2v��ehb��(�~�Yo�)5����  ��*ZO�����o�*�_y�+��W&���h)hp>lh[�;JY�T�X��q@�f�8d��a�謔0�!U�����5�(L/�Q��&=+�`�jG�p�9�F�ǎ�-u$qz<�5y]i0(�-=�t�G��S2P���.�Ǖ s�	�IF��Kׅ+�f��M4-j�<�&v��)Bb�H�G��}q%OWǱe����g����������2�sMKn3����Tv��	Q�ܳ�=w8^/����zԮT�yc.u�_*�r��}��J�94h���r熖$�3v�a&l4?�Ul���׏�S4�{��N;z�2ի�h��������M@ǐ]I�)�\�M�n
�؎`ш�& �{����l����?þ�C�b�5�����J�8a�8���LdS8�K
5>[��|��f�,} ���o��+Q^�'�D.HE�8`x��]m˙M�J!Zdj�Ã2߲�6�f� R�Ui�nʙ��\W�r IG�ba��1���զ�ʗ?%r�g۵]r�������`w�T��w��M����r�-N���י�z��h��z���I�����H�16,d%`+C�߀�iڎ~�=.����E�S�-!���ڹ��)?�Y�=֎I�}�����zg��f�Xg^�➧~�X�و�'H�! ��b�^�`4܇��F,P�Cf
�d8W�k�o�:\����.��F��+t1M�6+��t�+���PA�ï����d	:��c��г��3����a�k�;?�z�]ؙ���p4�[w���Je��M�*U��/(S���>)ڦ��5a�\d�ʙ�x_
㍶�M�|��,�C�zP
tݭ�ʣ�m)��ml��+�a��\��߷*l �8�R��lL��;C���M,�f��|6P�HSY�]��2+S��am9�Ⅱgx]��G����XV������\�����/�����`�AA�����D�"D:���*��4�#Hex�U]�.��rF�����%j��"�7���xL+_�&,ͷ�[����x�6���:O�˙z�ǯ���,C~�u��i�8R��.[,��gw�+̡eRA1�Z�������׬����͆EqJ���p��]Q��6V�Z�|�a�$�\�F���1e-������I��_?(� Y[z|���C���<�k��9��1Q��y��i\8[�m8\�S�'W �����8_h�cM�r[��d笟E�31$�J�\�.)��q'y��M4�s���������"�h�*�f� 9�F���8c�J��58�qpB��3��u��[,�A���Vh#���
8m�H"/�
��p�l�d�a�����B���!M֘V��fl�yy$$y�TInD�������)S����,���X=�oF0�?��ya�i����R��~1�Uy��'^� ��SR�Ax)�H��,�T�Ĉ�3>ظ3'���p]]PJ��N�d��B'�2���������l5��DP2�?�OWxB����Q�"M�X��ω��P�q�����8�P��7���L�7.ˀ���k����j1�E3��q�aSs�'"55�EgW�'�%��|����|0��w�b�L��9}�ߝo 𞘳կ����*��\>ԩ	jU-���f�:�Q�8�(CS~�G�kLo��vKԖ���g�[���vhS���T���!����]q9vH�2#x?X��ئg�iLD�z�X��բɃR�$&a���G].�f��P=K�N}�G������k����8���gj�۴�ǲ����&܎�����Wxvc�?�3lyn<1Ez.
uƯn����aǹD��nv���B�iE�� =<Ę��u䘄�'rŉ��� *�D�{���C���Ţ!�?,�Y\xOt�fF�"z�JD�mdh�3}n#+�
����C����U& !�����n�� n�\Ϊ�O����V�\~5�-+h�0_vы��*x�&Fؘ�q>��(�n��f�2�$�c�mZ٣�U�J6���L:l	.c߇TZ#����Wy�0�[Q��fjӞ����l��������V~+o�R�͆�^�Wq,~��� {��x���Q"J:u��K�FON���;�h{�o����י9��G6OuFa㾩�=y��a4�*#��X����v��,@�d�����b��&�jpM��?D�*�e�o����$���F��_4�p��A�#^Ǣ���&B=�<6sb��2z�/�+��MP�R�`�2D�r��ƔB�A���v3U[����w�Q���ђ.�LA�ă�3U=��p��"���[�OLSmh�ղ�r�tJ��	���꿋P��E�t$�_W� .��Hmb�IW3�wl÷�S����k��l���������?�Dk�(��l|���7��J�-��I�Ç$LB��ڣ�_�b�o��`�]�"��>RM1J$�{7��J�/�G�*�kf�Щ'7g�d �zC|�ˈ`��;�b���Z���!m�%��Y��>�!94`ӂ��~6��d��k1Ax��Yi���=�Y���e(�o��S���2)"d[����(��%