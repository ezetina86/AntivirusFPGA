XlxV38EB    14d1     611J	�-"����Jh��?N�V��^R�\�
�Jj���>�-�ٮ����v7�T$n���L%�R��n���X��'��y
G=��xم7	��b���_�����_kD��#��`��VX��B�G�:�R���$������BT|��C1vS��ܙT�� �"�Y��t��'/��k�Bm��$	eDIK���`3^%�@��-�L����?��T*0yۋ1CڪX�˘]��_����n�����DHx�j��V,�+[׭?���n
��h�������x�Ev~�S�Z��y��"|���So�8M-���@�'mdoTu -f(#��p�[���6��t���̖2|J�_ޓS��?+�����'q��X|\ت7M��c�U�Yuwi��4{�-△����8qu��G�E���1�R��:!9��JSV�&�?��G��.*Sa��\��i�������Gc�q���|(e����2�:{s���e.Ƈ(�ǅ`���/V�����5N#��TZ[C'����<T�.���. �`�����]C�uu�9U�U}3�Y���i�e�����4ݶB�s;2��i�9^��5�n�W��V��O&����ӡ��)�q\�Ul]�!b���yu�m[�cWĬ�Mta�g٨�^C��=� ,(���UjRZ�S�픣���Ymmw^���-�;���@���y~�J��Cܠ�>�Y�F{����f`��T"h��o���HTo"�۞�
uhw*�j��8��B�G&߿����[ɝ$'rj]��\�r�>@K�;�OZ��,���U��4�#�H��H���ӑq{җ[�#W�����e8c%^cu�����m~��ıb�js�4������*Ѳ)��z��:���A����� qi!w\(��d�A5&X�ж��v�=�Z%$���Jr�!��E��a{�+�r��RW�za�^��������υ$���C���#Yk> ��S��B���F%|�qZ=)]+��7�{:�����)�M-��/ߦ�b�!��N��ۖ��b�'j�{܋�g����r�H� x=��EV��;����P/&y�.k>�lH���i������y��e�itC��#4|Ox��&��3�"�mn:;�!.3���KG6��2��W����z�-���?��H�ZI�?�	���T�"MKW)xb���v�^�{$����= q�|H�C�i����%]X��D�f9��=;�I$�<�f�B j��i��`�?SMo^͝��Dp�]�]�*�<���YQ_,�$���Ћ_0�ۧ|6b���d���
���#%]�����d��y∝\;���n r�E��MF��W�E��/?}w��n�q1c�,�<����L����h�V�m,����g
!���uװ�FV�U�1#*Z��Y�u���]ܧ�KGz��3�s��Z�q7��ӟ~���w򸋼.[֊o������C4f'u��N@�wE�,��f�/�>0K�'Z��8���T�_���?�v'ó��#�zb�׸*��k