XlxV38EB    7c29    16e7ILL]�DI&�4�HM����	t��P�iL�l�؊�W�yo�0$��7,4��o{����>��� �s��'��	�d��F�ceK�&/!{�h�c�>V�䅌#�T������I�Th��ߩ��EpЮ��h<���C�R�H�j�b���!B`^�-�M�cG5�>�g���{�9a�u���8ORePA��d�+/W��<�tϨ��j�H9���qOc]�X�c����Z�r����{_Vy��H��~N��%UʢEܱX��ָԊ�l�$�� "�͇�*��s�B�Z3&V�y����J�Փ:5yiw����W���76����g��i���u��$�ba&��v�C�ё�_i�'e�T�����݀9l՟�*�Eav8����п�ye����9vc�OH`���-�᥈+M�#F ����#Oc$��[s8 s��gw���q|���o+�QIgb�w5Br��,����)Y�M�d��DtnX�J��9D��1Y�oS��u�	U��'V�MF�,x��q5[@���uW4ͣ�*(��,�M�ƚa�xe���ܶ��5�6l���V1��=`G������m�pJ2��>�i%K�6��%6� ���W�]��!3ѹ�0G~��[�����Ói_�E�gϵv��J
�1k��혵�M?M��q����9�$U��xHu1ǔ��
���\�d"_�s�����<,Y�bb�T^1Nx�_�^_`5:�(��Ɏh�
� �������t}���B�����n���qo�� �t�f-8��v2�:j���"_�-����YP�MK��@��i��+��խ�MrD0�s�yg�PD���(����]%8��#��PX*^�a�2`��N�P~^ �~V��=ܫ^�O�QVS�M8>�ʸ$�D�y\�["3�k�[�&]���B��h��W��9�th���l�/��h^t���c���q�M(��|w�Fy>g�3ݻ���c�F4��~u�dꕏN��9gY��Wy���{�R�f�x>6���g]s)-�8}�v�l�B�ӆ)�X�]]\��<���䴳�-7֑U���.-����<ׂc�������( ������<���
+"sM^df�lr{w���Y��|v[u8wYR�v3�^Ґ��ϙ<2�&@bh�'h�h�<�jm��1��S�4C=lT�o��TH0�4���;ϔX#�tj���g�邎���,�)��cc'��|~�g5��B�X�|kK!�k(�ً�F/��t�uv�jXӱ}��U�U�`��NsY��F*��/�S�j��u��z���D����V������w[�f_N�����%����ŔD#�k&K�7�k���	��e9:ne\(N�u��\�q��۳�J��%E�������D�����Y#�3JM��X4���0n�/#AZ��,G~]��n.����<�1p����z�w�� pz�X�Zy�aF]9�#��#��h�Ы�6ա&���4�MĢV�LQ"�ƒ�X��&d�V�ܝ�V����?��%B�,}�#Xq���������C	��8�	���x\T�М�֡{!����_	�?�XR{Eg�]�(m�蒟M�"�}!~��J�i�ǁ��ߢ��,�Ьl��������vU�-����.V%<�����Id��BD�ą���4�e�]�,W�-̢��z��lw�"�b��.������t��q!#��?M���e�,1K,��;�/�q�a���R����t�킴��$��n�_i��C�	H�"독��_�彻3޻~��kf	sS��s��v�<�����y����i��� 8���eq������	�H�K���EI��@.���m �$0l�&��ĵ�����Fg㉘0UR��ڲ#�=f�����!J?�#?�Ƃ������Qt;��	B��~Y98��K8��� �y����̼�34������_�*��l�����t��U;KQe�CTI�[�v�9a�w%��Q:�Є�މ�qs'��F�[�;�h^���~-^�}#�_�pj����$އ(m���zۤ��6���G�N}�ّ��J@�l	Z���BM��KKv�/�u�����@7�[e���!�iR��%������,g8'F���ځ�siC_N�!�l��M��/ZD��+��3|��n���a��v
IQl&�1�J���q�8t$F�Hb����G��=R���Z��f,��Y�]��i��wOL��i�"c�O�����M���^E�rg�����i+�?
���J:lX}[���NF��IF�0���4l|���R�!���2��D�m_��Ta���xk�؃D���B�?�4�wK�eL�q=jt�Ol���2�d|S��$(,B�o�HS�����-���U��f�":�a,+��rd��;T�P���-��\K�^�� 9!Q��NI�vI� R!m�)��>��/�T���Р7�.j'&ѩ��E����~?����g�h ���{�lo@˘����V$�=�&���h��nD�P�s�B�;z������ KZ�	]�`C{�9�/�[`z"{�$��o��� G����7\k�D�d;_	=W:�� A�@�J�&�����>q'?�0k�Yl"00xF>�����,4�l_E��?��)'���C�g�����	rm2�/��>�>[>8���S����9q�0�ax�Ig���0���٣}�/_��7%�  cb��v�z�H��y�lY�u7*�[`�`��N���i<��FF��8$���/_�5���N���pv4���-�*.'�^��a.:���v�CҒ�7�5�+�eô�['�솂5!�tR������An��sE�Z��s�)�`#U�D�U�mZ�T���%�]��唘������zl���ٍ��?���qz�O;J�	��p@�}Ds�c������
��<�$�b]����4Rõ����1��_�(v�pc%�۔�퉏���:"���G�L=%Z,���Ѻ��5�/��k�ڈ��5Ph�DR�1�K�$����o��w�F��}#���|����<�=�s׹p���)�kT���CKq�ĎDr�4��V�d��8eQ��H`���.&��ي>�<�l���O�}�6C#p�#�!ZzJ�job��8_\il��8�3��j��AdX�Lf�L3��,�uI��'�����
��$�{���4CB���2Ya+����5ټvN�5�g���; ������U@D��y�����a�4h��)H4�j���(	��v��#��G
� :� Y�Pr �d)�]����M掌LQ �3Z�� b��J��e�L_���uNm�@��2#�Q:��lI[��Y~���X�fʜ�QE��i��*��V�P��[����m*�1�]�ؚ4�3T��ŘB\���6#�<Y�K�A�(�(���0f�M�X����д�'2�O\*AB�I�S��T��v� ���v./�����P��l_�TK�@����i�jte���s���`�k*��[���B�vl�`^O�Y���ې���1��X�����<��Q�3a&
S4=h�A�?�ΖT�X8��#�����@�+�D��	iJ�z6� ���>`�\�H�u
1s�"^!��>��s����Z~��=Df�h����16�鹎�`����5�� �w�K����8�+�1����Bk����3lw�@m�*j~���I&�J,�i=�X������T˨ �wY\�ą�8^*VD?��
���#kq6x�� ���&�s<��ui8ZD=b�_�B�Ɉ��&�K��v^�,�{�:�H�}� �}�[�w�r��D3[�!G<����|�x�yM����˺���Q&�9A�gn��/p���w���>��$f	���-��/h���W���۹�iE69��O���*B�]���<F�GI��D���aNj���"k���I���G����i�GB���eF�8ׂP	���R���T,3����]Cu��(������V��W� ��TK�@gƳU�L�_���,�<NNv�d�]�t��g �mK��4J����;��i����+�.���I� 1t��J�G[�|�̯�8�ސ�"�DMj&7&�5���q��x�ܳ*��j�s��!b*����_��ԖE�#�	 U��H;�@9��i���e	z�R��R ӹU,�w���\�"y_�)@����O�P40�QK��>�c�2q��@;��:V*C�:T�z�����}�ZM�%�x�l���#�t�R5��{��Vn�Z	3=uX�}a��6�wo�~P��n/���k1�Z@�c���h�H�cI��T����qδW�QZ+�/�%�d8Nz%�'I9_^n��悒�}�*f�IZQL�=?������ �y��ص�2�ƣ�o`�QҷL�&8~�9\��;�Y�$y-]j�����l�r�{��6���l.����w�a�Vrj�T��%�f>�>�9r��{��V���dɏ��qh�/��Y�@��!��O�p')�`��K��Y��t���s�.�Ȋ[R��E:6�ָ.jz���.�RI6 �oہ�tO�[��8�X�嘓/�b�:�%!�X�褾��)�
`�Ň�cND�ө5\i
3=iU���]�J����*�G�b�K���g�C�B�)Yo ���c|
`���G����5#|�L�4&�i�H=�Дw�i�)�
ve�N_�DX���fT	-`�-"]MK.�\l�K�2+63�e��"'[�}����,�SJO6ci�n��㏟1�.�_��3���c�� �w�\��i�:�Ծy������FP����.d�~.WR���� �'$��ģ�Z����`��1���Db�E�N
�ֈq�����ci̦�*Y�e%Kܡt�7L�K5�4�;B:mPz
��o5U}wmM%����G��*}��-�p�ޏSLq�]�>O��M�]ߙx黗��n�/v"�`��&����#'Rs͖���S0.Y��9AQ���?Q�����u9|�\$wx��\KX�t��c>�;TG��õ
{31��O�������l�L�;|�=rh�����`u��[3fEj����Nb1|<��Yu��;�l"9�I�w�4�ͨs����s��dx�y����b�~�V��>�"�B�U�yH�]Xd���H��ԯ�p RG�̩��7��ۋY���궈�0���a?@o=
��;�
��]ZKq��{��sD���l�WS�\��}j���p�u��/�xV0Y��:���W� sf(̵��A�X9�HM�Ip���~��TW��\�#��~�Z!�/ǘ��"R�#�0�%jbl�Pص�*
�|��4�`��GQڦ��LM��L�H_N��*��jr�;������3ozf��O_�q\�)i��cWn������TQ52�r�o*b~�n���x��!\i�`�f������b�#��'�$���Lu��ɵ�أ�cw�p)�=�j���2�52��G�aA��.�!n��h\iL�-�{�`��׿�3$���x��Q��$e�,�)��vI���o(����s����!��T˧)2���L�s�	�m���ɥ�t<e�EQ<��6B$�����W~���L���b�2�5�#:�ZI+Tǁ�NP�oh,�~��e~k�r<��\Օ�{���s_e�8�YOG��F����X�!�i�jV
�	���ذ��$�kN V��e_I(����I1��|��=����O����l*���/�F��M;�_|�ܦu��cf}�hsP�W7g�\8^����