XlxV38EB    141e     4fb`P,�3���9���]
�K�bM�M�moL�6�5�*��4F��6;߳��%3."S�$5w����L"'��Od\F�*fcj�T��K�kK��a�&�cH6�a p{��p��_�u-h]V7ksby�����0�h��+�A�e#E�2�h�:���N��A��j�G[ 2��&���)��m���CAϷo��3G���3�M�1d��|2�!d�Q��Rm��/��#�ak4覹��f5�G�ȼ�u�����'o3V�hϤTc4�!I3e�<�*�jS;M��m�a�� ��G���c�z�q��k\�+&n�u��2^�ay8�o���q;�~���ܘ��^茂b�޲B1�n�J`󝀄��ڦ*�e��GqJ5�\GM������M���w[!m�fqz���sbZ��¥�^�
�.w�A�}Q���˝�B��U�����'؏n>1e �C��i��;BL�8|>}�+���v`b��IHi�,� ,"��rׁ��&�}y��Og3�6D��I�?_��L��s?�:
C����]�: �\9�ͨ�n�rQxc�
�Ǩo�(8TYv���HV�!�*:��މB���g9����I��Ƞ�9��K���J�Ѯ�ެM\��h�����_�&gG A�H����L��У��/�Uڐ�)���Tn
��a��8��O�A��83_��v�j���Ĥ#�%mj����o���*�D�NVC�oS�Xe���X��ٮ�1sM���F?�|���V�����`n�0%H���Y.���%
��aҁY.�Z(m��E��.�
�z6�MϿ�)�OW�I
./���J��{9e�ʐ��u�)<;��w�f铯h��%�H�ɵ4)���/z@(�Y)�ۘ�\^�x��r{��	�#�����v��K�� �'�sK�^F�O� �|)��	�>�(��l�y���U��\7o�9S�d�쿄��n������ �	�{<;
�1M��Gl!s6Wd�[j�\A0��F�)y��zb�s_�N�PW٣*/+�O�b���$��KqB�8��".B���F�G���ےb=d�D7�rf;z���2;�Բ���!��.� ��0O&'x�5�m@�:V4?V|*��X-�~��w�K3�`������=f�u˔6Z�H�N��WS�x�#�����\+�h�䇦����������ug����.�^�P� Ž���Ȯ�JT(Q�֖�cO�~/�쇋�I%���2Ԓ1M�?g;�R�����