XlxV38EB    11a4     4b0�6j�-{`%7j�ٺ;�^1�ʎI�0�w���E��C�~��<"�z��iA�X�A^��#�(`�L�l϶%~<.`��#��H�>��ۓJd��Z�2�������]�;@ݵL���o�cLU���{eF����g���M�{M���,��0���x�8�#�ഁ*~��{��1���~b�L�;� !�3z}m�L!�)b�&B�e���5di>5|y
Ȟ��a�:ʉ�EX� a�>1>�]��Š�0%�����2>d�X_�a�iݟ�N}��)�43�F�Q���.�R�E1���̢9P~x�I/��H/񗍾@e���L���?�,z��>*��8�ãD����U�VU46�?��E���5x��E ��?V=�A�g	y��R���D8�X�b_��	��
��\��{NuM`A�-�4$�vk0�5F?^d���T��->')+K����!��K�{n���d�8Ȕj7��{ER&� 3�!�l��Vs@=�F8oO����1E,#T/���W�K�D�����ߜ�J��h��v��K���G���� 4� ���jk�,5��;�,oZ*��}�u06Z���E�]kc��!���}8K�?ٿ��kI>U��2f��2�׭�҉8�t�4�E1͂с#, c�5����9<}����bruk������>{��]����0�z2�]�[<>�Ε��$� b��c��+�4|x�Q�����P�H� ,:y��$�^#�:\\3��&��	ty�J49Q�w�R���Z�>L��&H;T�,�"S��X��54MP���q�ܦEO'K��\À��ć�s^�א�Rs(�/i�	��������CI��"r;_-x����p`�)`�����p]{`���z#��v_�b�S(q��D8���ѫ=y"�_��lOd9	�:�F��_S��W�Ɂ���$�-���ޣ�X���a�C1ɀ���m�/��i�M��h�@�Þ8�?� �F4�ri6j�|P�)������0}�����%�R���|ƆҞK�+s��R=#*?���!=I������א!vsG�y���n\�A��J�d�nv�'���O�/�:��A���������M�S(�3������O��hf���[��K'm"}��}R��|��T���+���%:��,��9I��k��}�|;F