XlxV38EB    1331     4eb�)�C�y¿Ycq#`>!�{av��?x�j�EN�e�٥
��R����@�Y�N^ߡs��^JlV���d��4�$�1;7@��N�k��Jq=Q�r#JN�E�G�8�m��0;%�q�:����
�"�/��.KX(�M|Jw\�>R��$A^�㈾:�f�n["��1^ѭD���"���(5ך��ϙOi����������D�U٤��C0��^u���$��r���c1$x3�\�L���JYd�F�ϖSS�-&���w��D���zjSTD`x̂�l��J���0�����a�{��峺z�_���D3�]�����Q.E��#�˕�=�0o��CW�Pϲ<����6�w:oR.��/Jp�lA�^
�s��0�	�R�I���,��C�|��>�'�W�a^�tlSG�a�SC,��v\�x�6�U�"��s�� yهw�%�	����GIO6Yd&�z����UMU�L��V�P���1W|T|��+"
,o��A��y���B .���tδԩ��]>G�W}����Ǘ30M1��:�j�" n0�!��2���'	h}ZS�pY�69h��	�6������~�<q#�Vءy����[OF�w��Qio�S��c$.}	Q1m5��Ȝk�1�SV�D�6��ʚ�q/' �D�n����7�����zGg�Q9�q9R:1n�����ϋi�.�߉Xa+��8�O�adl�9��z�"�K�P�4�o���$xbm��b{��k��fe�<Ϲ�I��Q� Jю�sWH�����F���Wy��G3&3��
܄򭩐^�-y]���,�
Z�]�R���42&��[J�\e�/'�Li�[�P�ġ	T���o)���w �^A��A���T����6����Y�3���&&�Q���S,����_ "�Wdy�T[4�\?\��T����ה�\ C�"�ol��'�ҭ�"�#y�ss�N�٧{MG�P��aq�7bh+�B2Cv�����GsXU�{_Z�;��ʡA��'j?�T9��Y�[��b���5
�d�=8����ߎEH(���l.�����x���ˈ�g��9MаŤ�vte�ꀾ�9����:k��ɇT����*ں*~�O�g�҅c�.y��#D@��U�ŵJ��/s�quEL�z�2��l!�YgL�-bHp�^ƚ"�)}�@����8À�R�s������Hi:��;Ro/�Z}�jp�ܤN�u�T�J���W�}b�
