XlxV38EB    1389     4ff��k��Dt%>�¡]4Y� �I�����%�6�W�E�E�il;8�PL �B�G��Uk;�DS� �Ҝ\��\'�^���fk���U_}ͯ'r|Y��d��d��b#��.�r�<rC4,���c��U#G��G�������&�_�����H?��3"�A�������E-<h[м71U9F:$�*h�c@L�I�d.6�N'6߰�L�j4�9�%dNd.���͇���}o������&wDtrKһP=Y��kZ�+f�	�����u������O0��uwJ�D�q������`^�b�a�z�]�7	w��@�ô���l=�j�%���-Mc�S8�7����<Z���=�&��Q��2Mo- V�HK�U�^���1��@��C�5�
sF�����-5}��(<��B�¸��������El	6V�=nh����qMy���p��c���[�o��z��ؾ�F���*?e�������oH������i% ќ?��~\u�/Ϧ��%q0�
�.�4�S�2}CW�|y�
o�:qL�O���nXqëߓ�E�c�t{���0��J��� ��&e��]������W��:A������U�M�E�`��i:L*Ȱ���C� E�}y0��҇�|�54v}#��.+���zF�J�:�y�����3G�J2�p����zIIl�jd/�X׭ �fa<{���%�b�<6c�k]�{VO@p��7�<��Z���؀?�������#���^���|���C���ޘ���!-.����Fշ"j�y?��s�ގ4%-��_'��Єo�V��@����&��V���|��d
+D�	�[{f���7��PZh\���ZQ�V¨�éZ&1��ah�B�h	ī��\�wL�/� �,��
���]�W+A���v+�C�$���*	2n��]#��+-g{��w��+_N�'
��������@�*�,	͢� Q�%��`�����v[����1��5(�`ȣ|K���#�?��装V�s�W�ޓ뎅D�����.I��*�����`f��V�Dv	 ����)M_�񹇓@�0n�al�Rj���U���_�96_���ƨ�.1`�궳�W�\���{/�Tq��8�S _�iE��k��*u�fJ��-���r&�A��Z�l�nLjk�E@5졥���TV��z�яT�/�u.ݧJvԔ��6�;b��Q8�{&Uh
���3���� ʧ��