XlxV38EB    a946    1b8d��	�g2���DB%�H�g^��>�"���O�3R�B�%�U<����+}e��/{�R��m�3�����[���UZ?)�N�9��7d����*��2��
ߡ	�I�zF������Y�ĊI%��T�W.��*O�
@=�ј��w,�E���Tu�ŏa̕	��#���a�+h�7�]<�;���P �#C���9��������鯠'Dx��^���g���J�{4�����d_�G�=�ʱ��/zm��8�$����Oh\,K��E_����[����S��nK�\��ɾ�*�6��RqhT#Qa� \���1����R��hl�z�]�@p8=��c�Lnb��ԡA�o>����e TM��|�m.�$���͊�Ihőh
1 T�Rդ��0��J�>22VB�e㴸7P��%���Y.I�@?ZC����D����jb�f��1Y��CWȅ�w`��sU�@��05Bk��3qСz��G#H�;CT#P{�1�c�kv�P3e��
�|�5���OR�<cB$/+�ϧ�P���4� |3��g���}ny���61�+��⼍-J������tS�*����o7@���Jt�pAr���ꌓ��ǋ���$�T���I�p_Z�zjӋ��9d'�ԀwL����#ؤ���Tk�q��aR ��-s�~`\#�{}�(�Vg����U�ktӴ!g�>|x>a;���l=<$":>t<˔�is��̥뀮�P�a�'Ӟ�/yf�B��k�x��|s/#yM��O�ۤ�F?���2R�\c�T�	`g<t��1���R%v�S�W�h��F��J��Q��`���޴C�E��k��m��L���u�������PN��y)A�-t�K9 h��l\��^����v��(T(zQ��֗����s���iGl�ٯ���&cP����,G5�����v!͒į��Y\qF�q
%U�\����80���gS;�d3�����O?���3^Le�=����hg�Fy���v��e�G&w�LnWG�*��`B��]���ydB!��;�ԡ||��g�|��N�o��Y�:ֿ`3��4}��d�>^��j�n��l�њ>�����i��8��S��?d�*�Lt.�7�vIB���߂\���Կ`R<u��h
/ �M���\���]"�.��5�C 2?ḫ2��IH��=u��md�� 6#G�Wl��ٸE!���a�8���L���Ρ%�he;�^�慆s,��H+{t�‐5��#�#�������������/�ٟY�}K�j_�_s.V�o2XG�B�E�cة�ǅ���@�lM�ʈ��X�J�s�ާ�D!=!��߫O�K��aS2b�9lw�X�R��
	ޕ<�Q|{>�(�4�;H�W��P$���&� ��J��]m��\��=nS���Q��nuT��1���Z��v�B���jwm��U�x����U3 eq�9�SbX���rIeUE3P�G�
��Ĳ�<�}	�8ğ	Ղ�R��]��^X�!�.���#[Zfu�rf�;�B
�l���!5����h�����!�ieX��q'�e`��A�� p��3SR��������"���\��k��2r�jN���V[��@,��	�V��c�<1ښ�ݫ*��Dsr��,4K�::M���ޱL�0���;��΁g@��?U��K��a���jh0��8�e���E,n�v'}�4���l4!_�rB;�F�(P�s����7���Ai��c}*v(�1{܊���R�,�Ca���x����W�&��]���(�h<�05O��J �'��l6� ^�j� 6��25W{t�f�B��`��5��fA��N^�e\HD���'���m'�8Uc�P�a��r���/�G¸f�-,��dT.�D�_��°�����S9S��(��
8t��B����1(OA�����G��R���T`^,��t�@�0��g>;;�ڦĩN�i�"`è���NvtDR���[8�$��������4�6S��r/��v~8�X_�m#���u_a#LQRL|���P��[�{9�p~w�+#���79�(������z�*�ϴ�𔃜��)ȆmC�,+Ä�T��:��ͤ�(F�i�N6ǃ����7�T�⓼r�b��`W(��w���A�d��犲)�T��4 �;��5Ҵs�Q�)�"��i��	��pY���h�9��q@�p�n(ιr+ڋ^&~HB����#��(jt}��CR��,�K&��v̜\[�B����m��3�-�BT��_JxK��ka z8�f3 1�[p��9�����<n�,��י�&�W��O��8��˺˓���zD�����N:ֹ�7�B��m6MGK  ��]QD��$�/�?Y~�
��ul��f�KIќ���Ÿ��zUM0�%\�+5��_:6�
"�9�_��	��6�,�%_��m.`L&�X�ݠyx�#�2�v>k�ce�t��&��E�g,��/�	ٹ��|�l�W�n��H�����a�m0���͵el.oJ!�61@W� J����n@m32B���/mD��v�,BC������O�N`ȼa�/L��T݃�F(Q���33�Q�[c�r�k�E�Q�ߨ&p�{q������S5sM���ʜ��v�U��y5��Ӭ���4��֖Vq|n0��^kN	���>�A�]��c��|���TZ!""��Y5nD%�[[O��K��Zr��v�I��P�[cL�
3;K-t�*K:5yDЉ,��5p�G�(�e�N;�>ش�>e��;��+(�Z�ޘ���&��}}����l�_Pj��{�
6ޣ��������:!ɀ����q�Vq�MNŰn�(a�]���2W�3�)Y�؆�F���^-��،It�R�pE��<;S��:�����р��JxQ���KT���v��'d�
�I���V���'��A��,t*�"?�L�C����M����A\Tb��L����`)�?�����p��p$���s4��6��8/�J���f�yz��]+�(W�;p'���n���i�(;!��&���6A��*f��^4�.�s����U��"h�M�S>���ܟ�kˑ^�R����(}���:~����<1�׉J�g@��}zB� Q#�+N|�t&c�ɐ��s�qf�r�Z��#-�늎�j����*���t<����J���e���j�"0<4�@��1�N�U2} ���`E%q���z�MT���_7�z���:�Pu`�9�l��A�:9	Fy��"���L������&�wz���|�g�^HQn�8/Ԭ3T6�x.�?;B�Ϙ�w�W�M��ΙC��m�y�-��TZ
�v�m6� ����&�>��nܠ;!��������V��ʮS�W)#��F]p�u-t�Vu5�j���H�xX��	���ȡO���%o3��"ߊ��GZ����Ow�Z=�ez	1����x�0;���{)*��S�~T�7��y�%r���cm	�����$t��Nv��64�>����i��~{��l,}���ۈ. ^�j��&��p_5��SX!����(k��D��h��.	u��.샹W�4�R��߈�Qiw�m~b:0�?����>M�����u�.���E-�LA@�������dAE{<��d�t�E�/M�[��P�4�>ߏ5��t�<
@ִ�S�l�:$	�- �pe	|lQ�+�+�>x�6%��.��Ym�C�.>\C�b�#\�ʄ	u�8�����h1w���s�ף�t��˾�z�neh�N����� �]L�A,4��� o� �
�z���p�^Ư}gET|Ø�G�W�P*�x�Т� Fh�	MÄ�$���N��Z�r�Uz��$n�?1�vaO�ָXӰ�S�X_�䪹ց��[6���H�	� D);d�Ox��c:�-V��*/2:c���{K�E(IQ����H_ѧ���Ƙ(�GJv�{��Ğ-��Μ�mt�OPpY�(;T���p�����t>f�[�:O`��su�i�z-2�{�e��������	�VA\�o� ��(ǓO)t���E�_r�EK]&�1ߊ�'��E��t�r.C�H})Q��am�nFp���0������ķ�2�E}O�ܠ�P�]Gn�흨��>ɕC����3�#?�D�F�w�W�����\��W,���+�!��$Ť�ĘC@6�H��:șWBif$i�9���.�����ˆ0KL�Uj�FO���"����>
�Y�q���3�FeM�Wyg;�p�����O�ox��<��I��#�s�N��ED�{R����ӼV�	�<^�=6~���h�Z�B>�*|~��Se9��%�G�?u�O���??r)�D`��P!r���"�t@ �.����R-BGa#�����`�n�E!�Q2��3�<{�x�pN�^�8?\T��P��<���*D�sœ��s�Ȭ��AP=��픬vB���)�y\����5z_��*����? H~Я6���+�>ʨ|���N��	`Sn�����o�Uu�`����#�#��Q0�ц��a��z3E�"���'W#L2>j�a��o=a� -+qa�� �F�[����h+a��t��I<�r�X� ��ņY���H�tS�X
Z�����f�q4�S~n�>n�Rq�����v\<"v>����3\�q"�|ֈ�9���b��w������ H7/M�(�;4������&�v�ŉ6&��f���@LB�����:�j�A*�4�>�/�8Y(�e��l���P[j̆]��C&��uӋ����l$�o����R#7%O�Ay�����z����pj�>�*�ĭ����f(��@|9p[�*�^ȏDZ�E���*s��޻N�dC�	}�1��P�'�\|g��^�G8c� ��i��#}9�Z)%�t*��/��u��6�~W׮���t�6i�)�q�1���c�?J�B�ln� �����'�2[�}SÁ��s�O~��h�Ճ�2ڬ1��q����Î��b�Gb���R����A�.�t G>R��q6�3��_M>��;F?lV�� ,$i�����
��V��~�C�1�f�62����K�C����%\�0�j��Ϗ�|�� pB��̢�u�ש�D��M�3�Us�J'��3`A���\�qt�q�]D�z}9�?�B5�G�nU����8=K���PO@��x)��e�͊�o3�r�)R�`[�=��}��ɮ1�Q��}�ww��Vյ_����mM��l~��)6
%���)�*,�`rp���\,�H�_@;k������}��B;P�h�K�9Aƀ�}��c`�x��3��`�"�H���/6���n,�Aν�2��D��Pmg:e������xj�]x^}�e<Ky% �Ug����ɿ��&��O왶G_���xDAcߣ�=�#I�v�,��R����Ƙ�|���u��C�����S�;�����H��n-o���{#�1p�H�b�#��e����|Oj)}9_���/�t�皱4X^�!�Z��:B��%[��!�p	p�G.ɀ���)gi�H�$=˅}�'�I	uF}�	��x�ԩ��la����6�i�cr���7Y?�(�G�e��Tہ��������aP>}"��6�M��Â�'E\���^��xTI�S򚠰�J��yOx��}ةyW�� ��bl��~�SzO�#���5]]�ގC����C,n �w������Df��-e
Z	���8S�� ���%jHsY"-y=��E��k��Q���o�u�bBHE������}Ez^��^q�#slTG���>G&s �|v�W�������k�n0����ƇP��k`D�����Q���& �x(�-1\��܊�>x9>i���~������r��U��87ߨn��������A����Sp�����v�I�{�&_�|��
,p���l��\��8|�k����;Y��݇jXQ��}��9� ��k�����P=��˅�j0ʗ4*�pL+�����|�"�0k�����v.l��
ˉ��n��c	�:i��Z�qC�-�y7<oVn�F=�"<����3\<-R&qf�xz��\I�g���Y8l�n��3�����U��kh�B1��q�Ի��2��pP����B;��5 :)�0b�6�*?�y;9���p�wݖ�q|�y%�?�{G���eM���:)�1R��M��)�}{�|Yخ��Q�Of���_LH�����TY'}��y���a�~��k�(��K�̊���x�;�?Yg�~���7�,�U��M3n�k�i��f�Fl��������+򇿙��6�.�Q;��)saz�+��N�-vL	["s%�~B�k�3`�"|��m�QT��4�8�,�)o	F9(S�P� �cs48n��yn���%Elj��i��!��
�ݾ�yɃ�K��������X�l:��>P\����F�l]��NX�l�����"�����IF����_Ү��A�&��r���Z"_��~/�w<�;	���r��!2,7S���6na�UZ´��*2W�ު}\�[rN��~y���nhA���Z���ٶ��-��F����# oh�Et�m��B��fN��j�"yecs�X��9M6��bo�3�`Rߘ~8����7+l���k�D9��A�����Q�3Ο��|��B��!7��J�<���#�X'�e���u��S�J��|�=�,o���R�N�r���&*��[bǀ"y����0�K�Vm�����m��sAe=nD�d�u��f�Ӿ���|� _�l��/����3i퓘y-q��1}�d9M>�=E��}`��J�:�L��`��N�F�p���v�/������0E_,@���mBB6}YCS3 ��9q�3�Q�n��d��k'�l+ZH�͵d�����ݹ�|*auȽ/.�L