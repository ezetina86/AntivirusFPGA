XlxV38EB    146c     52b�#�ꓳFv�����u��܊��0f_V]͝�9���6�[�eBa��N{����3Tg�ڠ��G)�8���Փ�^'�\����!�|��ɚQ��l.��jk�P��t��g�]�g()��~,t0�&��<����X��[��<��Q�ɍ��P��.��Ȗ�(�$>�v�]��
r^uďS׭=�\�� ���ji>��>��l4��-��q�:a�)ăɵ���9�-���޼Y�v���
M�ʻ��֌v9��w����5�`}B�`w� �13��m*�u�Q�rʯ IͨI���m��^��M�p͙���\-�_�Ւ��pIû�f��Jln�u'������1̦w��Пs�LCVF�?��	��rYY!�����ɛ�~�bb��y���'���Aq��YV�YC�e�%�I�}��U�S��lŴ�c%�\���(���Z�[�O �y=���Y��0F���c�)3-h) E+A��߲��a�:ݕ6��e����k���7�k�ӄ�-P��R/� ���䒄�{��%e�a�w�.n0r��&�
�7eFR�Mȴ�t�w����*`��1J ���jZ��Pu��5;C�as燾`[7��,�6�&`J;�����߻�O�����D&71�S�ig���6��wܓe��NF{��,@?+�o�]����ɢ�\��ç �0H�zD���;�e�5>�ﰐw0����-��A��+�y��CZ	��MHag�%;�"��^
`�~˹x��/<�]�Ȫ�_� ��]~��������&M�vm.%�lm~8�5�hJ���y�'Q<>6uY�D҄�o���O!�y������0%�~
h����L3j�NnJϯMa�iA��B���=�9�U'�l��t[�,�����3F�s�g�[$+HƋI\�6�W Q궯ȗw�� ڡoĐ�@/�Ҥ����qCT�Zo����@N��"��k�w�T�+��Gq	�+UM��0��bs�Hħ��g�Ɔ��g�Tco�!��Q�n(hcN�,0�"�}$�E�����̦hg�3���d��Ka� q.V<�+�[>���g��1`�����T�q�D/�AI�>-2�%�1�������xx&�+g�A���I3���&<�̐j��wܗ�θ!�3KG9�3ר�4���0{�-+��;�)}_g-N���u;�2lN>��}���][h��s힚I�K�Kt����E���1���'s����tU
�,�����86`��R"=onn��
u:}�G" �A�D����~�X����,�;�?w9yd8c���2Q��l����X�%m`R�