XlxV38EB    208e     a2fpW�]��..(<��^Y�(zW V�c�%�F����x?�l�i��Hx��u���R5\�f�LH��ŏ�q9M�
�p
��;m#XB�!&Y����?���T��1�@-(�o�pQk��P�"m����g2n��A@";|��n9��n��P����s�e��(���+�Y�X��5��H\S����"u�oK�!��V71���9FDb0�fѷ%It0�B�{�X*_�ņ��w�w��ĮP�@D��5#��jj��?\��'H>c�/��I*�87�w�����s�u���݂��$����`w0���,�c2M^l6w�i:k�f*~��F�Z�0���-=`�FxD�c�jÔ)G�!�U��Ĵ5�)��Of�@���S������~��Q8�Jl��X^WF>�]�Pp�msȱ�w�k�K�O�iD>�����P�>�D1�>(d��o[kg
c����Ƿ�Nt$��M/�Μ�te0��ل�_X-�{]C~׈�!�Z�Cv��W�H�*���s��m����Y��t�#� ���p��	�"f���cm�ln��i��9�="�/�nF����C��(�7���{tʲ��H������$���{��A��T���)��W'�U�_���������h�pFn3
��IPi�2��O	n�`���'r /�rq�q�hl���:����B�Ca/bI�H���փ.�u:̿�����p����Ɂ`�x�xŝG*1[s�EXG����fB�8�3͐��.���a޴��*���W���&_m�態p�Z�y�J�J���F���QW6�A;.z"z�9ϯ#h��G��;E�8��ȉ
5̔�����
��UR0?��b��^?5�
0m�fm�й�"/d�r״ϥ����o�Rt�R��w�{d>ZD�Aq$���N�k�à�T)vV�x����+��k�N\�[_���^ӷw*�\ɗ�_���f��*^1� _����˔�a�u���=㚽~�j���H�<��� ld<����ΏN�`.�Y�Fi��N��N��샄 H�L^uiy0���u�����6�l>���������Hԉn��5]��������3�a�z��3i����Ҵ/_�������4j��0"�����s[$�rZ��4[`���cE��1����Gg.����W������mo�?�<���:/&��U>�L}��/�"���܂7�-O�PD�{SY��D���{����^.O�;;�m����ń�tf�L���.J��c�(z����/@�ǵ*�)ϊ��v�+>��;U6�(�#��XU�z�Q�9�\`�ix���SY|r�"���M�}f��x:�XN��4�r��X���֑I|�����#)o0��L�u�aE���f�v����mXv��@�6��Cv��\l�o����j�{�<�!��2�'����I�������:�o%�Y^���Y}M�u��ͱxYA���yl����kg���ȏ��.A����jrqbŮ\�L�,�ϪS�5�Op_��ج��������w�GɈL�5����4��%4�[��&4A��=~\�	��'f�i�m���Yg�.��E� @����K�S��%J�0r�ը�;h����A�d'T�x�(��EZ0����o.��l��߅s@�1�nN��B���0n��A@v�y��ȥ0>��z^�\�`�PI'Ks=�Ƨ^��1�
Y�ȮJ.��\���D8�7��`��v:e�Rk��GKN�(���� �U���V��A�f^5t��W2Im&�iG� ��:�ΏQ�%�ڋW�\�O!
ج����`^e��CC�Ye��X�>���T�	�<���~��VG��UT�]$0� I��)�<��u��Sw"�-��@���)&W��|�H�g�*��8��<�?���<2�[���o꛿Qz�y7���؏ �Q`���򜓝�UwCe����Q8��1ri��)�V��O��]��P��΃5LH?���5���պ.Y7��rX$�2�ז'w��5l�%�`үE�ǒ�$���e9�W֎�0F{A�~NxUq"���������]I�ty`'���YI�#C=I���+��c��!� ?�ǯ�.�$j�~�xU$D�������#?�R�{3&�%ݥ^�`��NKDxSP8X���k����;9b����r
�đ"#�h����9Nb�����m<&�a5�*�}T��#I�O�~�_E֢�ӆ�x��W]lt8�Ϧ�'����D����n���n�vR��ݢ� s
�6�N���5CE0��g��́01��~<�Y(	�|��_�C]G���u�nv�B�"%��Օ�Hq����CZLMX6hR���n�M��tf�4�^�$��f�a(�T| ]�4A���闑L�$A�_���z7u[w��*Cf�N{��� �)s<��YcW�jȒ*�J�J����WM �:�*�c��j�Zs"x�/6�Q��?Hg}v���a�ߡf��9p>f£�\�-Iԭ�vE�ĝlc���j�T���]M�hV�ܼ;�1i���T$/pg���
�\�ƌk��[e