XlxV38EB    1442     4ffzH�H;��g� ��$��16�j@���Xj�ܠ�K�9^��8�3<����ގ��"��NkK��B1F�M@�Og����z)rOA$�o�8�q�00�_VR�n���)����U��F�1����va�ZY��W0E����)$bOZ�[����+:7�U�I��qV��]�;��$�x/u�o
rǼ�b#�M�!��eן��i(ͩ�X�=৾��qJtA�f� _/U�Ù���ǉf���GG[i��0C�g�_M������Xc� ��z	�;]�B\#b�0P��~9��m*P�Z�DY1�]'O}������!=���M��1r�o[�j����ɹ;E�z�<3s������>���]-�VCx&H:+;9u�:����ǖ!;�_ w�}�k�r����?	J��VR7*�q*4�Vq��mJְ%�H#by�L�N�b�a����rn�4������̧�eG�4���)��5���T��j�	3�`��7�����)�)���sR��Qgf���A�������C9�13不ᭃ�������ĖÛ�)6ڟ��z�^௲fN�|F��!i�ѵ�8��g5�V�E�!]�]�� z���C���93�y+��*�Zf����X}U��Ge���I�ͮbu� ��^�U� �ߓ��~1��+���.b��W3�9�=�~H	��h���0x�2cm��_:�����w��h� E~-���G�T����w��E�6�{-�ABT��.pm�Qֻ�S���YǤ��� f�-�^D�L���������6��|�<�BN:�Җ��Hs;[c������zI|�Fr�'���|�M��]0�=<�u����t %P��M��1�L�����ښfI������l�O���r�ٳ�1r;���fX�kl�1�#lɣxN���|k^"�ܼu"�zA}nD��6h%.]:���@L[.�����&p��k�G���Q���Y.vmJf
�`Y�~
 `G�*��z��u��Ϡ�nK�G;�����p�Xįv`���6�,�p�c)���*�(���6��J�r78�T3��4RM<-h���$i���si���T�q�>�%��O�F�s�+�2���f]}���C�q�ܩTȧ������x�V�`M6&1I��R�P:�K�7=A�DDc�/݆71�0�E��Y�Fms
�M�ŎY�_��j����Si���2��j��!_&��:6ܹyÙtȦK��zGsAWmY]�\0������