XlxV38EB    1914     649&+���������q͈(5*C���&^b����)yoNgS2W����;����~�~��2�K��[�oB��iT�������1��*�W6�⒦)5��z`
���"l���,��;��>t&�(&�������e&�$;�Ogx$����\�+�rCV��X��qiǥ%a�0�,{�%�a�{nO�c�=
4����ea̤K�J2�㪼d+�_������i�Q�N?M�>���v-�a?�U�����R��M�� �CB�&�,���ܡ���c��F	CK]N�����{�%+�w����xeK�K�vāݣC�]������!8[˝x[l=�y\�-c�m#G˽�Kd({�5�<��|���x��Hϊ����R�t��W�}#�(L�W��:��S���5��U��T��a�] ~�h�D6��Ia��4�oH�a|pG�g^2�R�v驗xH�NXV$�*���	���+�!*�N�g�X[\���7NLG��%�OdL��1ٵ�����l�.NA]'[����	�ػ���G,�um�"���L��1ƛ�*�xQ�}/^J�ڒ�4�ќu%i��9m�l�q`y�8�n�]�d��y(���0k&��:�X����,�;|��(�G/�b�Ѡ���+ *����Ԟ�B6Kh�����~�Rz�e�6D��*���t\7���b�oG��Mx�bH�^ʛH�n�� ���#�泄w�g=�Z�@8ճĈL͏bG�P����.p*��I�^=n�U��7�^��ͱ�����149��
���+��
�F������ "�No�y��R�6 ^���r��âC�o�Q�x��]m���Xb�v�T�y���-Hì�7$s�
��\^7��E_μN칉1#�	5��׿c3O�ct�u*��fI���F���� =]���խ�7D~�|�$~�W�A)
xC
/YD2���	����D/P�0��x��P�`w�C�sJ���R*U/v<I=�3�v�Pq<;����I6��������?2L�.n\�h��1bѫ#6Oaq;eT�:__*B��*�(�'7�o���OSt��? hL2^�A.C�7�	q��x�rdr~r�7�Y`#1�T�������0r7Y:@��/�5��������f4���P^�^��T.�DIC1��=�I0�%����|o!�0��v�b�6Xۊ�
��Iɳ_�>{J|^�U7CW��؎n>�o�z!˓��1}8��8 7�p�O��5�	� ���
e������+9� �t�W|P���(_<�҃ɶ4әXN� w�F�i��~e��л���357�0Sa���B��2Qe�l]���KT�z�l��8�4? ����ĕ)�_���o��(lI!��K�	.���©[�U7��e���>��p�L�>ީ��Sϕ�Y\�)�2 ��8Μ��X�
ZNu���]Ǣ����U�w/1��2��S��OA{NG�X�}��̞Fܧ�E��Vז5��ؤ����|��Ǒ���k�d�I�%1ޡ1�(��D�ً��C=��c�tM;��)�Z�-��n#\�bcҺ�Ջ֐��x�T���T����