XlxV38EB    11cd     4a8�)�C�y¿ɧ((b��=��޴����E*�f(Cfs f����Ǘ$,�̓��r�=�����AGTԦ�R��D�Pv��:�P�����κ}�h=�?���t�h����,?ZM�Kp�P�:VJ+(ڙ���R�/ѧ�d,����i�f�a��@g��I����9& �*h\�-/v�e�U���-
�ޤ4�i��ѳ���~�8��kZz.IY�X}.G��]��<uw��s���~r,jn����7��FM�9KI���tό�˹:��=�x�̶6g��%��!%[h�����	��'2�+y%K%r��t���݈Yjw���ܚ�'�K��;��u�@S��4iC�}�	��n��O�0䭭m��y��#�e��h&:/���>�S���Rҵ����b�D�' ��**9�*t[Y�	gE���J�9�3�-��w0E`NIq�'f_9�������/��H�Ϲ��\g��e"MH��%rtX>:����)!I [G����nv�a��ΐIW�.r��c�M��z_B�1H���N�@AzS�n7����H&C�	�5VmK1��n���������J�} 6��[~�֣s��sz/cR\�CI�����D��M���3B���gi�%Ą��Q���r��|�a�"=�3�UF�cҏZ�7Q�*�S������dj��˭�"ph�q�>����Q�ef�/��q�o��"���xjt@�R�%�d�SŲ�S�{��o�t��:y���-��F`��ޙpk�\��e�\ $O�	����J|f��HP�c]m��kz,�w �z=`��1s����D_}�8P��A
���h&�|�����B��TH��W���kLB�������aݥ��Ee�Xc�j�[`"rr�±YgO�?饿��&5��<���J�r���
 @�hT#�ipa�5���SSa`��LA�R���߇ޝTН�z�whsom��
��QD�!3ޝ#ȭD�"�Rh&���rp�Q>ҙ;ߍ����&�OyGe+�ytUK���q`mH,���Hr�*3����փ�"K��u��;T�T'|��(M^@�)�cGi&�@���D��v|N`�#^�"B��o٧h\S��[܎~;`-��*���Oq	���2��x/�*+� �r����x��E	O[��!���57MFQ�