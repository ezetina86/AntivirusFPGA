XlxV38EB    3632     bcek��D� o��7�(�^V�ڙB^E�;�b)���e���ϰ�0J��Ȁ�kIxp��Rr�Qd����p���S&&����=��e1��&���[�C,����0�!�w�>,�/x���� E|�!�Љœ%�Y[��~Y�>ʞͻ��w�z+�%2��f�V@�������;�/��L��e]�Ywq��z�^&+��M2/7I�_��2'%ޜ��Q�X����&�"B����Z��J��O��Wx�z���`���jQ{(��e��@�΄�CE���HP�X4:��)�D�٤˴�)�ͨVA|��1~N�(>@&"��3��\�$U&�)Უ^���������aS7��m4��o�<�-HJ���,I<H=�~J�����Uu��]�S����|�!�O(�l�0E�=|�R{�o�[K��e"�h��� |�]��򐄐Aqz��ܲ|Vn/�0(&�^������$%�����������?DbZ D�j��Й��2�UhT���<����9�M}f&�h���t�'n���� C?]��e�z�/#L�%|�M��$WAلĕ;���|��N�#�zodo`�'�e�*B�1"�]�{!��J�@R�+I8��ߠ��l�;��ͦ��� ��C*J6��$���ݤeY � WO��:�B�iJQڤs�~
��α�u���D�a���]���U�^4{ާ�������G5|���	F��Z�~k.��D�\�� �y�Ŷ��[�q����� ��L(>MN�O$�[����UF���%x(ߑ��^ǹe�xz�x���3O�
`4#��۵�ۈB��5�V2S��[�p~�.Uf)�� %�P��;��%-$Um<=�)Sd����1d*�P�{��<7�>�l٦b�(�ӟ�����l4ޙ�|���ء��i�֭�gm��d��	k/��������_Te��@�nO��S)8̷^�����0^+�z[k��p�oP�'_�����Q!z.�H�3����(g��x��*Hj�/�����?:~'QH���⬈|Й$�9�	����-iK�?<�b�
�l<��w7�T|�`�6�Hy�}ڒHa���	�e�G��y�~M-�`%�E�~� _A���|#�k<��(:�[|۠>���& ���M����E��ە` ��E��s�l�#��tХ��� V�`.nh;5�����cy4\/T��5����=��K�9�t�!�����y�v���])}�͖n��gk���,��V�U*-��sK74��?E?C"����"UC���3����M��B���X�k��@.g��K,�*���v��ʕM�JVW�����"��S���Ғ������x(�d�}�!Q���w��`{����i�Y��c]��Nj�9ѡg&�c*nD;���i	�v��c�g�3��s8��}㕦���o�?�1�Ѽ��jg>�q��Qx�Q����ݺ>���)6��i��ʄ�a'��my�R�>�ӂ<��N�uS6��1�"��'/x�4�k�G�94c:� Yz���ҟr>J��AH����nnsx�����Ƃ����˗�A����OrĜ�r�`1#�����6s­V?�C	d�Ժ�&Ɩ�~�Y��3S6�xZ�� )����%8ަf�k���C��F��4���2)��aPo5y���'Ѻ�L�6<ME����� $C�����e�aP� �����=�z(%^!�Oż
BP@�l�Ԟ��Z������$PIq搼i�0'�=92�p�Q��`�������Q�+������; U
8"Kf��������U�~��K�De :���嫾o�(��#Cȟ7V�2·�TI�8D�w�K/�t�x<᡻d�2�I�0\EuV�=�@����>|�|�*�Y�iIS���69,Ǉ��}��q"���aV0s$���ı՝㨞(���rm	��a��������e> Q�̰�s�10�R�����3�o��TPo1]JLxc�Ay�rM� �D�}[�Lh���nFo�!<�`�DQ3�����-�Q�#u�`{��8�����vjгb�+z?���e�< �w'���#�d���o��w*D����U���S��4a��������	�i�o����.�O��Ffi;'�8>?r{<�/1��
O��g�R�[���oD����~Y��_u��CB1�����}��������>���C�H�������r}��d����x%���Z/�d��w�(�.+qм��̛]	��~��/��^�����C��a�y�'"��J��r���wqm���x��V�5��W�ĉM�l�z�;J���M I8j�2��b.���g���6�y�����w���a�m a��\!,]�^q�NJp�W��]�����Uq /u�IE�2��x.�MxŴ��� �����h>F�^�찷��E����/��H|E��%�_� O������t/�9c��k���S3ŝ3�"=��`X���'Ö�ۓGk��	(������|
��4�e��9h3�U�y��d:��x�������l���t�7�hD���1⤼
���^�Xފv9=z��	!�%�/�jp�l�XBJ5G���hBwU��|Hڏ�!��F,1��t郰��񥊁�Y�-�T��ӂZ�����_h��h[q��I&�,����ָ��jm�P("(���>1k5�_��l	�[�:�N>��Gn�4M�ӑ��{����
|�21��5���ϻ~��������N/�o����I�}�$U�W��H��?m���Z/J�_������R���,��^�u�"�Xq탓���R��R*��ԁ����A��i<q�&h���r9��^���ri�K'3tXO��7��++9��:�du�&0��_9L8����H%:��f��.wS/���1�I/��Uގ�:�X7S�m*���-�*�����n�zc�G�+Xצ
���?�C�