XlxV38EB     4f6     19e�e`���tFUU�c�m�t#K��D"c#�	ECSiNW�$��8��Vw7���t^����}�Kw��>i��������j,�d�8��\z�i���gm�1L=\�������ֻ3���m�1R[ƻv�$r�v�OLz �g�Z�D4�1K���#b�_���=H\�Y\�k,O�|���D�I=��LB&�#��k\�tл󙵸�[c�_ ������A��5��eQi9^q�7���]i7}�:��"O�ݒY����~����F���m����o�C�Fɳ�{ ��%q�$j�Z�V���m����V�.�Ta�aQ�2�r�QB�q+6�[��@�s�?�XHx��"uY����֐i�=~��hS]�j|j7IE��`M �j|���f�:��a���Я���mO�5�?	c�