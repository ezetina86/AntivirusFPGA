XlxV38EB    4d4f     edb�8L`�W[C4ym�'�Bi�y�Z�@騂?�u(���?��A�/�#���[x�n-
��'�� @����M�c������a�?�W�XOޔ����QJ.~!;��=R��-�m>6a�CM�ܿ��n�qnփ꼸/�����ԥ�Q}�$W��?�i�e�6Ͽh�֧��� ��!��a�K�R]e'B� aMG�s�#Z�1��������7 ��}8\��!�[U����#F�,-�jGD�B��>�{��S�̷՜����|����i����W�*s��U/�큿�j����D�8�t�
;��h&%D{��JD���Մ�9�$�f�ɖ�������>^`�����IQZ~!���:��V���s�>�#�0?�P��ܕ���'8�Y��bHd?)�G���}�(A���~+iej����gߧ�ӻ��$A・�ʋ03"��R���4ZU����28]�/|�i2�]�
��h� ��F��0]��.`5�����Mm�3���>�Lg�f �{6��F�N�{�{,%O����� Gez�r]��qou���9�FK���eu�s�bV�.b�-(�z�����4�cf�y:�ZJp�!��(٠A�/e��L����_r?j�߃���,Ĥ����ij��;��#�!	���DWk��[�R�I�']�(�юfV:�X������-�7�4�м���,J�I����g�������Z.zo��W�����֞�i:OۆD�q�4Ӽ���_61C�R���1~g�����N���IdnC�Y�w�W06�{���fx|'�dXN�K��X�7�~�7�iHB�Ʀ��|}��X϶/���	�q��a�'�E��XN���잌�;��"��^��br�|$>3ʬQ��zA�sh�j*3͗a8||
�j�_�R�^}�¹u/��:%��p��1�h�A�eQ&gG��4?WP/dқvJL��v�uZTV#W(�ϙd�L�k��g'���ϓ��[����.� ҭ�!�}�;i�:!p�A
��X��x�I�~l�d�JYN�	<W�Ni?�O�`{V,�HR��e��4��١�g��g�
�:�ׄ�0/+Q�xMw{i���ڌ:��[�����Aq�b��J3G���c�J/��D�&��V��)�w���<���	N_�Sf٠�x9,�%ikr�}���h\W�4����k� �R�2�j��1���?�v�/'�o���0	Az��\�e��\`�4%��,l)�c��'��۫���F-�p�F�wr�Yt-*S�*�k,�ߴ��u�W�|��F���7�rGg�~���u9�p%�s��%?��v�q�,=�O��Z�S��h(m�����/���\���N�yb�!uQq���.9�t��0��i@�������逬^Ibk����[��7�6JT�ħ�~$�����Ep��	�o&�K�d��i��n����|H&��Ιg�q@�w�:?��~`>��¿zR�7{G)ݟ��O��L������{#AO�R��
��$���7�.�|����`P��`(����>�J�shV�"�����ב^HUy�/ߺ��6���$R��"��B�8M��b�:��?݂�<鰷_$����h�v��|I�z\5I�f�_׌i�k�OIɨ���ued���9>�L��n_������mz�I�M�2�pV:o�]���ݷRk�_��k�B��!��o�DDg��$��e.S�δ�CP([�#@MX���¬���w��~�}�����u�l>��o[���B�k��!�_����=c�n
u?�j_�#�D��~g��r.��0N�,�&2��,�3�
�'n@��@m(�MxE^�/ 5H%���L���KR��;]�nOb񓺢[�xG�P�^�K�gE�d��j�����o�k�~��7n�]|�Om%������ �?�|On�H�32ǽMC�a1Dj'B��ҕ{��k����@m��;2Ҡ��l2��ֻ�~�T+��so-R�h�����-��=s��/���̃�I|��Q�$씇Q�nJ+��V�P�KR/�X��(�C����/����wH�c�:{������V4z�E�[m��2�j�*XR�~y���:�S���5�O[��^�{4�����Y
JQ7B�C��F6��:�ZI�m��c���劚C�[Տ���6B��Tˬ"QϺWxښ��Kj�Gj&d��t?;�A�#�/�M�� K�&�"A�$Φ�t����I�m���e�W�n^k���+8���� s��~[�>8�u��f�g��$�-�!������pσ��4��(n�¡aMuE��(���1"g�'h�Q���l�XU.�9�F<��ė!�z`%�B� �����q�֧B�\k�4+�Ã(2a�p�M���>�2pɰ����9������ٜ?�WO)y��[�[kX��w����1�2�(�M��} �]G
��c�=�P�ϯ�I&�-�m�[w]�"�����3��f�76
W�&�隃��H��-�~o1�����˜-���*V���cK])C�X�s�J�����"����y�F��ǖ�	Y]�:v�㍽�;<��oHh����J2����ql��S�����'�n'/3�sB�y�g*v���Z����9!lT�K�>����pD�Dc^�(�	x�/օ���q9�_�Č/����KebqPm��f�����mZ�4t��1�L��'�i�jO���/S���o�)�m#S덶!���nD���!�_Aje�.���:_H��43x�(��"�8�y��x�w"0��>�C�h�˩'Z�~M�(��OV:q���9F��z�x���sF��u
;n���(�J<~���5g1��P�,�7��&��-��|^k�E�zB�\$���ښ�A��ſ��EF��c����I0Pך��2Af���������&@�W���A��:�_w����/�3\+5}`�g��xD���Lu�sU�B�����}?	,�����]g-^Ȱ�2ʸPd_��Vd?j?�E���x*󐁤ܔq+�=�H�8��C�:&��p%o���F/�g�|����5�Db�lh�(�I��y��Ws��-X��V|��I"�˔j�%����p���=�HYʹ���V ڗ�C��#5i��J�.��!��i<c�+ܰ�r�yvo��#���T�e��!���]rY��F�.�a�pml�$
KxMe>mgWw�:K���O3��U��g+����SD�^�i�Ux��F��1�{e����I��w�y��I�, N��&L��yk6��N�)�Ȃ��p�7%���.ۼ�ͩ%��^p��ƅ	#G�N�����w0��Z���Rܪ��_CO����q7ړM�lh ��<S i��q�#s�<)R57�� ��c	�]��z؉L2��#bNJ��OA��L��S�DF{v[��FR[�����6O;
����#WI4��|�(�����q/0n�,-���������4V��'�Y6p4G��(~e"e�Yc��g9�;e/��m�
��1�_�����$�제=�g��ؑ�ˋg��c`�j�N!�8d����Xꏮtm0����c�s�*L�4�eOh �*A�����0�zbqW[|�S��{���%Gn���643w��8`�ｮ3�ܕ8y�֑H�'�My������qu�Eg�l&���ɀ��-U�^p�