XlxV38EB    46ea     c5c�3�N��)�L��TE1Kz`���}e�����q*����t�l:X#\��X���)���Ъ ?pZ���-�f]r��$d#U�)i��5���t*�ˤ��L�'��Ѐ�SQ6�o��L(.X���M��o���0Q8��.��76DG�r��$.O�^�L��H��C��c�n��`(׭���qP�Z��k�Y��blS����*��;'�O�X��v�)�o���U�����Y6�F�N��4PR%q�5nVQ:�� "�ߣ	
M��>��.���'w�V�y>fD�5�u��όmSn����n]�N�]6Z��S�"��U��(mU�HOz?̉̖��$_���^�"K]'�o߱�َ��-E9�ٜG|����a�J5�C��M_Qg3�� {8�Q��]::�&T�ml�F�Rp)�@�#���\.��H���Q�3e<�Y[('�t�s��U�v��H�s�9��Gm�ot8�O}�a�΋��}�ƈ���60I8[�P.� �'� �B�:���%)�%�Unu��L��B_i�����)��U���b
�3�
8�A`>�QT�@�6��V��SmѬ����9�DN��FO�d���5������p��||ʷ�����%"@
0..��*�Թ����X�wUgȸk��+���+�{贓�2����ew.��ά(0N� ��TX���=��>fVg��=X����^��o%z��eU����k��'����
7�s��=�"d4�����:��O�E�j����E�K �GZ���ޝڨ��/���A������.����]D�1����1�����n��6�GD��YA���X�����~s`��I��`5��<V�*�\�$&�J�E���w�kkp?.��TXv7�f�[�mqT{^���X�$b���c/��hA�IrA�Dź��%�)y�om��������'P��c�X�;Pj��|�����+�+A��c���^�9���,aWA�Wk���8&�A)�x�g������(����5Yڏyn���Qx+puB�i�qrsg��>��c�Mj��wYh��]y�� ���w����>��-�UD��OcT�����+z#_D󤕳F8�.|$�|52vCE+^�|E��5�t�­/�^'1>��FQT�z�si2�W��~�6��"` ~����ɂf��su[rP������#���Έ�o&\o�c�r�����cF|o�~��̍#��g&�SWkd-����`1�hfJ�K��n��νG�R��O΢�*�G�	4xA)ӂ�D\T�R0������O��k�W�
w|?D6Z'�'�}��t��T��H�⻑@�	@��ۢ4�_S)�^��+-�F�~d�z�J�F��p�y�rds�s��M,p4o�}���S:s�|��*w��KE{w�� �Kҹ�E�����2�^8a~��eՖ���د�5�*"d�ė��xj�������[7o�&e< �E7�˦i��)�>��S�mQe3?��<(�>8C����;<��ZFl���"���7�c?�1v����%�O�y�b���ǫ���V�A����}�qR�����ð��V� �ݹ␸�J,�29�v�vI^>�v���؞�6�� mڼ�Z)���/kҍ��C��P?�Ԁ��[9j~�c;*����8��C�C�'�|�N��jK6(sgφ�^����f���ު%	)w
hO���.�W	�,Y�)WaD�WuJN�m��k�c���iP���e���'#f��	�[��RVa�m�T�O��Lp�E�(�(�b\����C������!�.��x�]��h�[&/B�˝6{ �i�gu��� ��+띜-�~�L��Q�r��+ZY���W��$P�!݁ԃ�o�UJ�y�c�j^�>���|�1B3 X�X�75Ota�ދMsO�R͌�^Pe�ھm$&Z7������EwޚF�N��M���i>�c�̘0�N�Jw�	O�hkUs�Bn%.{���.=��+Ζ�8����Z�+}�1�[}a��Q�+��*��S��,�j�?��C��t�1u��S�(��r����e'n�B�6\������L�ѱ����v{˪>Z��?��Z�5TrL��k���Q����Mbf�*74l�[��ϱ�Ftڋ<�;Zb�<#s�+��8����H��|�z�z0@�����L�����s������Rі�7�S�s_���>q��**r��(ďw�:Kb�5;y^��c���Z,�=i�5�E�@.��P�'�Ӭ����ԆiIHb���r��Q0����r4�#��o��h�������#���T���:)=�
m�[�n}T�L�Q�{�2S}��9fԙ������)��9<"�pRw�?�˻�����L����Q[���<��6��?��{g�?�|R'�.>n|�r��vH˖��EJO�,_�J�a�>_������^m�mN���ZU��C��� �4��EJ|Ɣ�53;r�`ih�&H�5�Bڏ⊜F(e�-�nC�_�#��~bj�y�4ogy�B˱��b��ljf#u�1�����8ԛ����� �v�3�g��.��E�ed��)�}�z��!YꝖ �BQ��� Ev��f"sp3{�����PD��h8���}N�8J�Q�g��&�C��xQ$���P�. js��^����!�[O�[�c��Q;�(�O�O�1�m����a�4@�_|��F=��ۛ=z�U�ǃ��5�P�;�ǈvE\�����P\����KE��(b�FZ��N��Gk��_%�b��ZW}L�+d�E�,��ET�]��B��-���π�+C��@V�$'��~K���x� �eXS0S�-[j�'����d�'���@�ԡȠl��Y&�w��?%o�u�V�\��-�A��� eb�Ȟ�>0�<�T*5����,�0����D-E}1B_��������VC�7��t)�!>Kl�f-�H����[�f5����Ԏ<����2��r�	⍗�g�>�?Yx��wG�/����Yw@��>����j�E��Å��y�n-�F��#�7�Ig�珞��W5��ܢ�t@���wõ�k7�����~��q�fӀn���Bq�����!�W���m�e�?g�u��