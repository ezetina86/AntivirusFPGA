XlxV38EB    1122     471<�/��B�t@� �]�x��^&)�ҺW�q��8�H>�}۔�����1�?����T��ݾ��7Mw~�>a|Y�݇�7RzL���Sۜ�%�8�#$���'��|�v�V��q�Q��s�MO�o�wjٵD��_�'
Z�f��s�C����� ��Ƒ�׹I·U��%G�<� � ��ld��oeonM\'��� �_����g[���yDs+%��~J9��(3MY����9�$���^)Ӥ%7��%����&5@�*Ƈ{BAyE0t%A%�_�?������Y��;@/c�Y~0�6� ��xOD���srP<�.QX @n�w#�������B����z?�k�]{�",��G�eSrkFZ�X����P֪=N�
���%�5�!Ђ��DI)�����/$���&���z��C��1|4��g�����0���[��%�ޛђ�=]�i8/x� v��8�Ώ�	�M)��>�Ĵ����Z�c8h�7��(���j��������}�o�f`�c��DXFKn�b.{��Nx#4j1$zy��ꁓi��o�A҈��n�1�1�3�� �|�#ѿF��)��9 �����F�`X�s���R��T~��Yx�6�c��d��\�q�ZǦ��?�Jɠr ��a�$#jు�f�Llj�_Se?�{"�C����V����̈́X��m���$�#�	�ι&��^A�& @�8gR�;�D��RXötu��y��Y��?�: �}�]f'=�s6(CS0����f7)�S�7���x4s�܁(?=�㹴�7c��{��TD5�m��q�ˇѨ���I�3[�~�J0a&l�p�F����O�K ��-��8EȄV�R(���v�K�p�]�'+/:w���V
��W�}�����! A(������(ٵ7RV%X^�1�3�!`I��@H ��?a�-o^X
�1�n�8"���gF
s�i���<,�q��[��P'�ͣ8�$Z���b�1��'  -�����G�|��˰�n=�,��;�.��E�8&�W�-,a��¿]��M~l����_�I#q�
�=��j��%�h���Q��W7���wT֛�ab��5��&��^�(vy��S��k������