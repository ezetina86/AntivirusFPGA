XlxV38EB    1316     4be�Uɔ�Ґ
zr�0�	&�G�	O��VqLH������+�c;�Vu��&[u�'�V#����gs�h��B�c)2Z���~���nM�jN��̓��o:�X��pi����c�>w"���ȃú��x"�5uoԛ�����6�������A��sáT^5~Qd(�l�QD��&��Ҍhxtr��]'M( �*��3���GԘ��l��whx�\Ou�,!��%�uj=s\Z���O���B�|B,c ~-���Ȟl�A? ���8F��IA�(fe����O�f�q'���T�<���[zis�H��H�[��b8�Y��3s���jlE,_��ܱ+f���,W'
���MP��7Úu^)4��n�&����:���cg7A��+��j�L��y�xfጽ�����ε��{�q���=�PHN]F�����6�}2r�:^�>^$��Gy�{֐}B��Nj7�I��>��M��<���W��3.4�o��>kS��;Y��AA����gn��	[�`.��̈́3X�
q�]8Л/KIǋ�M��7�;�>;��𾉆颷Y�����k��e}��[5�����"�Z��;���ј$�R�M��آɕ,��*�ZЖ��~�����N��2��2�$�N�>��$�)-�֬	�/���v�|�n�s�h�^�S����^H�m���0s�Q�S�; ���C�C��[A���pzMۚ�����ELyi��%(�� �㭟;��i��Y�ᖩ���(�hp��]�X|�j�tK���b�x���)�����g.��9?^;G���Yn�^�X�]k���Y���F��*��T�W�YA����򾭙����j[z��2���#ƥ��(O������M$^?�&�b��f��ȺȫĐ<%�Q�hf�ڏ-xA1!��Yq马���F��@��8��-���m����:5���c��[3���P�C�2z��5���BD�M;q����N�Hf���`+�y�K�N�P@0_�¯i}�����]��MV��� �.ڤ�8 ��F�9ukx�ښV�Q���g�P3��j�y*�c��,Gpb>|�ǫ�L�1��Ak�P;�P�J/��Ky���)�#7�+�[������X%������	����l���l�HLD�h��R�ޚP0�:}yQ.Ó^n\��6J׋�?3q