XlxV38EB    261a     8df����fx�i�C|Y�K��F#ln�5�Ǯm.:۹�v2�LsGE���$�z�� ��F��`��	O�5�9(�B�=����5v�)��b/P������Q3	�TqM�q�[�'�Dԝ#��)��}k]��V(2"m��� ��G���v=�0a��:
��N�kJɒ�l��>{iC^����Z��mf�"�u�Ż?@:��uR�Y���{���[��B�<~n�q�HVceF�a����Δ#��`a��M�D�Y�0���j�q��X�Ia��q�>���ڻ1�~��P�����d-�S��r�����I�F!���,�wX�]lo~Ux�+�6���s�h�^F��4�.��2� ɾ<��c2�:3af��!�LCݡ�I�E �a���uږ�FL/#���e��|����� �z��k0��0�����܋�)Y�0��{���_��R����dΈ��ώ�&ҩ�y{���=���������fe��L��`�twu@�恈�����O��)%�3�]SŎ[��*t��`�¯�;�w��+�/}��t�8v*#��K?�*�����(XwSB���ˮ�2��������Zo�E@�Ǝ�"�o'+H�N�朕�TzN�S�;t(K��Hp����y��9����*K�ƀ4�t�
��4+ټ�����)|2����
psK�m���?"b{�v�p��8�羀	�!���!]��P��̚O��nw�вQB�o4��	��G�蛘�;�My�@J����TIƤ,�d�^2l�~�K����8��r��߬?�z�co&�!x״�b�#%s#��/���*Vt���E(_�P�����]{2k��\�Y�������8[hʮX��*~b�#����E��*�fS�a��l6���F���Sr���������8b��^�����/H�rNly�l��|������T¾�h���">e�$Z<�h*�.�<�+���n�;�mB>ܠ�.N)�$�d#�:W�>��a~*hMB��&���鍶`hI��3�iȠ4�����,g�
�Ȗ�?M��S�Y�s4��}��Q�����/ˆ�%��=�� J!� -3����*1PZNxb��0��Ǫ�:�z���R�aQ���̥t�J����d����>EyK�t��L��:bw��"�9͌�d/�9'B<��,�<o���F���R�ֵmK
b�N��9�wû�Y����aZyu�~@׍�Һ���O��S3�hC[*��<�,�M��=RG"?�&�ۓ�j?�P5'���pexr��X�1�k� ���48��(vmp?���zԺn�ﯢ4�q��+�z7,��x�G �t*����:=����"#�O\ePjr�j���x��༶+'wmE�ڣ���P[�~��t�FCh	��6L �^�C����p#��1����$��g����f��.��m��a�����fS�#���X���I�Nl�a�kEK�(���uCv���ܱm�8���Ӈn�\9�i�o���P���?֧���b�2�?KK� ӮE!�YV��[k�
�1x��:l�we
-@V=��)�E[�
�}.��l��|��л�0�����:#"�JJ'����Z��<uV���	|���k��#p�W�i���~�� �ɐ�io����o�B�3Q;R�SGI�q�K�㗫�ֲkHe���y���`7��`6��Z�����yޅ)8��ւ,�w7��#�x*����RK| �Ot׋T�rkb
�vfty$�SU�J]�P�E�!3���A�O�c4�-WsM˞�Y�T��p��z�.w)�#FNZ,�F��_��ɩs��F�w��[{9���Q�?e����L��3;i���C��#64����Osw�iy2��.��j�a��&
���qa��ȭS����9>"0��vYb�n�F�7�y5�{%ͦ�qs�U�N�|(,����`�Wo��ðE|u�
��hu�g���i�����Z@<0�} ��	 �ɸY}M.����mxN:�����g�G^���24b*�`W���~B�0�����S�є'�Z(�{o��*�%�����ٻ�P��C�Ig��x�!=���|��Q1�HfZ�$g���o(+g��,��*���Թ[���::�
��W�W�ӕ�=Sv��||��_YL<,�=��R���TeZ&��B��>���׃�u���8ϋњ�k���O!a��������D�V>� \-�h*�w��