XlxV38EB    3591     a66�����A�I����~����S�%��P:��;�܊a��Ƒ�V��K���%:���T"�`�6��¸���z�}DH���~*�e��úzB�2]�u�D��oz>gd4?��D*I���W����:��5�Ϝ�:�4M���_�Fv�DJG'_�u@��z	�J+�"�%��W|H�77��B`	�#�_F��E��:G1k�V� "�� ό�m�-:D4oC���s��K"E3i�����AN#��st:o۷ō����J�kӋ�B�S���'R�lr� bؒ���/�p�r|o �`����q{n�f�|dg@��ʶ���?��H~���`]������#� �5�Ci	#�p�pՁ�}v�Kz��Y$�+�Q��iL�&	�D�&�B �9���6#׫�.rsGX_�\�v���B"4�yҁߥ�d�gG%�%;@`�NJ��X�}�J��ǎ����p�czL�Ŀ��J�
�LD��C������z�~���F��5:(ㅓ/˹��e;h���T�SyP��?'k����Fh^����9�/�k����_.�猽��nK��+��k��%ͤ��h����Q��>X/>r�~��{��c�揮	���-��� � 5B0����x�I��\{_������F�%��"��5�P�M��z�yj���;%M�@�^�IR3�On���Z��S�v	����u�=�<�j�����/����y0%�<~�{�)L8��P�b�Y�u�q�8g�JR����������/�j�<�&���*�W���5�YNݸE�(c\T5֊�X���$�~��~ZGN[c��K׍>�&��n��?Ή������E������2Y]���k�����@ �k� ��q�[5�~X�#2%]�Oz���۪�j�w�`�}\�7&G�iO���5���8k\i��4�e�ŢT�j6�$����:��h�f99c*`^4��2�Yqբ갵)� �r4f���C�S�glZ�L��S�5�"E��Z��RM���`]�K�e$l^5O�>����A�|��]]��r�z��»>���Y�K~��uF!DQٙ�2�a?����Ý�0�5�bZ��p�����]���lSeǃbԻAt� �L������8N�� u�����I���gq�p9b�����ph�2fV��X­E�:tX����	�R+�%�\^��X��],!U\����$�3��E:��/��^%A�G��f;�[��C}�E�����p�@U�
�u7Y��d��`���Y�'ÛO��ɶ��/�`��7$����l��4�����J�;���(8����\�]��H�3�Rx%P� ��� ��0-�T�x��a�����}T�'O���< ��#RԱĭ���?Z�*)�`���J5G�޻��g��Lwr*�U;E��hF
���a���c�����(�V�\k��X=T��\����s��L�o�!���-��_ڌ>�EԪf$?V��3}�������=���ӑ���V��t$��@�N��H%~�5�+�|ߐ8�aUJ=,�O��̗"��a[B��D`�`p�'>�� ��"I�F���W��xPμSo�{�Y~��3�A~X�N-��Et:�(�Q���m�}����I���p$yb��0/x,�����_�hΖ)��������x���M��x
6�a}�#��V˥S#�g-�<��Ƣ�l�����M/��s�%�s{�PY#�r��P�m�c%9�e�e�p���!=��#�e	j�[����ݮC��"_�u�J�z�ρ�8�ݪ��]׏t�����x�A����=?E���]/����s���0����E�I�Қ�@B�K�&�5YA%�h/Tl0m����M

��W+�Bc��1�\�����[��\�����Ѷf~�pw���?�G�Im;�L�v�^��e��#f]���H�exI�{�wmg��(�� *��]�h���I�}q�a��$������!�.����k��G{MZ{���b	t�|~���ݷ�
L9������3A`�Qrc#˹{���݉p�%;OT�4�?ʶ�����m.$ծ�D��E�H�>�D�حZf������(��/|�HE��I�(��j#�Z~��xTw�CY���7��wK�y���f��8��偪UjBJhn���DHUn*;;�p����n*��To�N� U��xS��8���%'!�kh�?�M��X
w\�Rsob*�^z#��0��aW��R��4DT��a�%�z���u٘��&(d�
�M��,)ɤ�����x�9��JP>6��в���U9����7Z�m,��%��9}��n]�q7҇2��2@�O	/}X}���'b��1d�|�2;/�n�>`�M�
��٘��YR���=��INO������Et��XJ`n1iz�&,S����G�Oߪ�D)��J65��X:��,8��}s�E�j�U�umj0�w&�t4�[.}�BQ��>�wHJ�w��7{n�D�d��Q8;�`ys�~c�#�T��gD�-e��3`��V�a3+^���LN��R���y��d'��B�$�24����=�