XlxV38EB    12d0     4c1#H� ����eEq��I�C��Ӏ�G-7;f T=��еB(8Y����Ղے��O�?�m)qO�$���vJ���� ~�f�P�r!D�ͳ1�'a��2�$L=�j�v�9i^?=/&��MK�^s�rW��3���7�GZ��}��9;�_�I���nE�vV/�sb�Ω5>��L�?������%����Ze��2='g۪�*��`�G%�wg/(�����/��oE�IP���u6	>{A` MOk�����b9���רdl�}	VIٻ��!����7:j9M�\�t�uU/��vA�}�����Ъn)����^.�hn#9v|x\oʚD�cU|�<q���l��"�A�y/0��g��h��h���:�����Eֶ�1p���'z~sN��F�\!��9ls�1�b��:�Ƭ��yU ��X���F��[4G�ȃ*�;�.**���X��j
zxk�Е���e�R�u��?�K��r���>���+� ��g`�rp�L�q��%t�	��x�X38p�<���W9=��Kg�E��
�b`-4�q�������� ���������\����kݨ�6��K0i�G���u�dtv&�]HH�P!x�ɸw57�Dlm&����c��7�ʹ�Y�:$�(Ӽ�w{m�,Hw����)9�x��م/��9���O�a�{g��8�֢��!���������I?o���i��k*{'ބT�89n�&E�����dw▤�N���<���b��)����.�����q#K�v�Lծ�U���д5w�a�;�g+��,+M��V�o`��'�LhXd�F
p�d-I�,S�D���%��������1I޺=��)�?ޠ�gp���t.���V}mj�n��|���F�w�X�r����b/��ʐ/���	 "�d��<��D	\�3���.��z��;�Kj�~=]0�	�LX֓Qm1��HOuaM<?�h"��үݥS��l�	b<B�9Jܛ׎dT^eG����טk�{tF�����*��nU�S�m��\�eyO0p�'JC�JG�&�vh��K�}r`r@^N3`3�ԅ��Q�V�	�%O��D�ON��8$����z%����~��T��A;�!��	�j��GPǟ��[^��X��0����(#O�A�͇_�q�5�����`~��%�r�M�#�ɽиm��UӢ��qE^��E@�2ae�<�9�#vh"E��c�W